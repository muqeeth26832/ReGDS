.SUBCKT XOR2 A B Y VDD GND
M1 net1 B GND GND nmos w=1u l=1u 
M2 net2 A GND GND nmos w=1u l=1u 
M3 Y net3 GND GND nmos w=1u l=1u
M4 net3 B net4 GND nmos w=1u l=1u 
M5 net3 net1 net2 GND nmos w=1u l=1u 
M6 net4 net2 GND GND nmos w=1u l=1u 
M7 net3 net1 net5 VDD pmos w=2u l=1u
M8 net1 B VDD VDD pmos w=2u l=1u
M9 net2 B net3 VDD pmos w=2u l=1u
M10 net2 A VDD VDD pmos w=2u l=1u
M11 Y net3 VDD VDD pmos w=2u l=1u
M12 net5 net2 VDD VDD pmos w=2u l=1u
.ENDS

.SUBCKT AND2X1 A B VDD VSS Y 
Mmn2 Y n0 VSS VSS g45n1svt M=1 L=45n W=260n 
Mmn0 net127 B VSS VSS g45n1svt M=1 L=45n W=145n 
Mmn1 n0 A net127 VSS g45n1svt M=1 L=45n W=145n 
Mmp1 n0 B VDD VDD g45p1svt M=1 L=45n W=215n 
Mmp0 n0 A VDD VDD g45p1svt M=1 L=45n W=215n 
Mmp2 Y n0 VDD VDD g45p1svt M=1 L=45n W=390n 
.ENDS

.SUBCKT INVX1 A VDD VSS Y 
Mmp0 Y A VDD VDD g45p1svt M=1 L=45n W=390n 
Mmn0 Y A VSS VSS g45n1svt M=1 L=45n W=260n 
.ENDS

.SUBCKT NOR2X1 A B VDD VSS Y 
Mmn1 Y B VSS VSS g45n1svt M=1 L=45n W=260n 
Mmn0 Y A VSS VSS g45n1svt M=1 L=45n W=260n 
Mmp1 Y B net41 VDD g45p1svt M=1 L=45n W=390n 
Mmp0 net41 A VDD VDD g45p1svt M=1 L=45n W=390n 
.ENDS

.SUBCKT OR2X1 A B VDD VSS Y 
Mmn2 Y n0 VSS VSS g45n1svt M=1 L=45n W=260n 
Mmn0 n0 A VSS VSS g45n1svt M=1 L=45n W=145n 
Mmn1 n0 B VSS VSS g45n1svt M=1 L=45n W=145n 
Mmp1 n0 B n1 VDD g45p1svt M=1 L=45n W=215n 
Mmp2 Y n0 VDD VDD g45p1svt M=1 L=45n W=390n 
Mmp0 n1 A VDD VDD g45p1svt M=1 L=45n W=215n 
.ENDS

.SUBCKT NAND2X1 A B VDD VSS Y 
Mmn1 Y B n0 VSS g45n1svt M=1 L=45n W=260n 
Mmn0 n0 A VSS VSS g45n1svt M=1 L=45n W=260n 
Mmp1 Y B VDD VDD g45p1svt M=1 L=45n W=390n 
Mmp0 Y A VDD VDD g45p1svt M=1 L=45n W=390n 
.ENDS

.SUBCKT c432 N1 N4 N8 N11 N14 N17 N21 N24 N27 N30 N34 N37 N40 N43 N47 N50 N53 N56 N60 N63 N66 N69 N73 N76 N79 N82 N86 N89 N92 N95 N99 N102 N105 N108 N112 N115 N223 N329 N370 N421 N430 N431 N432 VDD VSS 
XU179 n178 n179 VDD VSS N432 NAND2X1 
XU180 n180 n181 VDD VSS n179 NAND2X1 
XU181 n182 n183 VDD VSS n180 NAND2X1 
XU182 n184 n185 VDD VSS n183 OR2X1 
XU183 n186 n187 VDD VSS n182 NOR2X1 
XU184 n188 n189 VDD VSS n187 NOR2X1 
XU185 n190 n191 VDD VSS n186 NOR2X1 
XU186 n192 n193 VDD VSS n190 NOR2X1 
XU187 N329 n194 VDD VSS n192 NOR2X1 
XU188 n195 n196 VDD VSS N431 NAND2X1 
XU189 n197 n198 VDD VSS n196 NAND2X1 
XU190 n185 n199 VDD VSS n197 NOR2X1 
XU191 n200 n201 VDD VSS n195 NOR2X1 
XU192 n202 n203 VDD VSS N421 NOR2X1 
XU193 n204 n205 VDD VSS n203 NOR2X1 
XU194 n206 n189 VDD VSS n205 NAND2X1 
XU195 n207 n208 VDD VSS n189 NAND2X1 
XU196 n209 n210 VDD VSS n207 NOR2X1 
XU197 n211 n212 VDD VSS n210 NOR2X1 
XU198 n213 n214 VDD VSS n209 NOR2X1 
XU199 n198 VDD VSS n206 INVX1 
XU200 n184 n215 VDD VSS n198 NAND2X1 
XU201 n188 VDD VSS n215 INVX1 
XU202 n216 n217 VDD VSS n188 NOR2X1 
XU203 n218 n219 VDD VSS n216 OR2X1 
XU204 n211 n220 VDD VSS n219 NOR2X1 
XU205 N329 N86 VDD VSS n218 AND2X1 
XU206 n221 n222 VDD VSS n184 NAND2X1 
XU207 n223 n224 VDD VSS n221 NOR2X1 
XU208 N370 N79 VDD VSS n224 AND2X1 
XU209 n213 n225 VDD VSS n223 NOR2X1 
XU210 N430 N108 VDD VSS n204 OR2X1 
XU211 n226 n227 VDD VSS N430 NAND2X1 
XU212 n185 n200 VDD VSS n227 NOR2X1 
XU213 n178 VDD VSS n200 INVX1 
XU214 n228 n229 VDD VSS n178 NAND2X1 
XU215 n230 n231 VDD VSS n228 NOR2X1 
XU216 N370 N27 VDD VSS n231 AND2X1 
XU217 n213 n232 VDD VSS n230 NOR2X1 
XU218 n233 n234 VDD VSS n185 AND2X1 
XU219 n235 n236 VDD VSS n233 NOR2X1 
XU220 n213 n237 VDD VSS n236 NOR2X1 
XU221 N370 N66 VDD VSS n235 AND2X1 
XU222 n201 n199 VDD VSS n226 NOR2X1 
XU223 n238 n239 VDD VSS n199 AND2X1 
XU224 n240 n191 VDD VSS n238 NOR2X1 
XU225 n211 n241 VDD VSS n191 NOR2X1 
XU226 N53 VDD VSS n241 INVX1 
XU227 N370 VDD VSS n211 INVX1 
XU228 N329 N47 VDD VSS n240 AND2X1 
XU229 n181 VDD VSS n201 INVX1 
XU230 n242 n243 VDD VSS n181 NAND2X1 
XU231 n244 n245 VDD VSS n243 NOR2X1 
XU232 N329 N34 VDD VSS n245 AND2X1 
XU233 n246 n247 VDD VSS n242 NOR2X1 
XU234 N370 N40 VDD VSS n246 AND2X1 
XU235 n248 n249 VDD VSS n202 NOR2X1 
XU236 N4 n250 VDD VSS n249 NAND2X1 
XU237 N14 N370 VDD VSS n250 NAND2X1 
XU238 n251 n252 VDD VSS n248 NAND2X1 
XU239 N8 N329 VDD VSS n251 NAND2X1 
XU240 n253 n254 VDD VSS N370 NAND2X1 
XU241 n255 n256 VDD VSS n254 NOR2X1 
XU242 n257 n258 VDD VSS n256 NAND2X1 
XU243 n259 n260 VDD VSS n258 NAND2X1 
XU244 n261 VDD VSS n260 INVX1 
XU245 N115 n262 VDD VSS n259 NOR2X1 
XU246 n263 n213 VDD VSS n262 NOR2X1 
XU247 n264 n239 VDD VSS n257 NAND2X1 
XU248 n194 VDD VSS n239 INVX1 
XU249 N53 n265 VDD VSS n264 NOR2X1 
XU250 n193 n213 VDD VSS n265 NOR2X1 
XU251 n266 n267 VDD VSS n255 NAND2X1 
XU252 n268 n269 VDD VSS n267 NAND2X1 
XU253 N14 n270 VDD VSS n269 NOR2X1 
XU254 n271 n272 VDD VSS n268 NOR2X1 
XU255 N329 N8 VDD VSS n271 AND2X1 
XU256 n273 n274 VDD VSS n266 NOR2X1 
XU257 n217 n275 VDD VSS n274 NOR2X1 
XU258 n276 n220 VDD VSS n275 NAND2X1 
XU259 N92 VDD VSS n220 INVX1 
XU260 n213 n277 VDD VSS n276 OR2X1 
XU261 n278 n279 VDD VSS n273 NOR2X1 
XU262 n280 n212 VDD VSS n279 NAND2X1 
XU263 N105 VDD VSS n212 INVX1 
XU264 N329 n281 VDD VSS n280 NAND2X1 
XU265 n282 n283 VDD VSS n253 NOR2X1 
XU266 n284 n285 VDD VSS n283 NAND2X1 
XU267 n286 n287 VDD VSS n285 NAND2X1 
XU268 N27 n288 VDD VSS n287 NOR2X1 
XU269 n289 N329 VDD VSS n288 AND2X1 
XU270 n290 n291 VDD VSS n286 NOR2X1 
XU271 N17 VDD VSS n291 INVX1 
XU272 n292 n293 VDD VSS n290 NOR2X1 
XU273 n294 n295 VDD VSS n284 NAND2X1 
XU274 N40 n244 VDD VSS n295 NOR2X1 
XU275 n296 n247 VDD VSS n294 NOR2X1 
XU276 n297 N329 VDD VSS n296 AND2X1 
XU277 n298 n299 VDD VSS n282 NAND2X1 
XU278 n300 n222 VDD VSS n299 NAND2X1 
XU279 N79 n301 VDD VSS n300 NOR2X1 
XU280 n302 n213 VDD VSS n301 NOR2X1 
XU281 N329 VDD VSS n213 INVX1 
XU282 n303 n234 VDD VSS n298 NAND2X1 
XU283 N66 n304 VDD VSS n303 NOR2X1 
XU284 n305 N329 VDD VSS n304 AND2X1 
XU285 n306 n307 VDD VSS N329 NAND2X1 
XU286 n308 n309 VDD VSS n307 NOR2X1 
XU287 n289 n281 VDD VSS n309 NAND2X1 
XU288 n208 n214 VDD VSS n281 NAND2X1 
XU289 N99 VDD VSS n214 INVX1 
XU290 n278 VDD VSS n208 INVX1 
XU291 N95 n310 VDD VSS n278 NAND2X1 
XU292 N89 N223 VDD VSS n310 NAND2X1 
XU293 n229 n232 VDD VSS n289 NAND2X1 
XU294 N21 VDD VSS n232 INVX1 
XU295 N17 n311 VDD VSS n229 AND2X1 
XU296 N11 N223 VDD VSS n311 NAND2X1 
XU297 n312 n313 VDD VSS n308 NAND2X1 
XU298 n263 VDD VSS n313 INVX1 
XU299 N112 n261 VDD VSS n263 NOR2X1 
XU300 N108 n314 VDD VSS n261 NAND2X1 
XU301 N102 N223 VDD VSS n314 NAND2X1 
XU302 n277 n302 VDD VSS n312 NOR2X1 
XU303 n222 n225 VDD VSS n302 AND2X1 
XU304 N73 VDD VSS n225 INVX1 
XU305 N69 n315 VDD VSS n222 AND2X1 
XU306 N63 N223 VDD VSS n315 NAND2X1 
XU307 n217 N86 VDD VSS n277 NOR2X1 
XU308 N82 n316 VDD VSS n217 NAND2X1 
XU309 N76 N223 VDD VSS n316 NAND2X1 
XU310 n317 n318 VDD VSS n306 NOR2X1 
XU311 n319 n320 VDD VSS n318 NAND2X1 
XU312 n193 VDD VSS n320 INVX1 
XU313 n194 N47 VDD VSS n193 NOR2X1 
XU314 N43 n321 VDD VSS n194 NAND2X1 
XU315 N37 N223 VDD VSS n321 NAND2X1 
XU316 n322 N4 VDD VSS n319 NAND2X1 
XU317 N8 n270 VDD VSS n322 NOR2X1 
XU318 n252 VDD VSS n270 INVX1 
XU319 N1 N223 VDD VSS n252 NAND2X1 
XU320 n305 n297 VDD VSS n317 NAND2X1 
XU321 n323 N30 VDD VSS n297 NAND2X1 
XU322 N34 n244 VDD VSS n323 NOR2X1 
XU323 n292 n324 VDD VSS n244 NOR2X1 
XU324 N223 VDD VSS n292 INVX1 
XU325 n234 n237 VDD VSS n305 NAND2X1 
XU326 N60 VDD VSS n237 INVX1 
XU327 N56 n325 VDD VSS n234 AND2X1 
XU328 N50 N223 VDD VSS n325 NAND2X1 
XU329 n326 n327 VDD VSS N223 NAND2X1 
XU330 n328 n329 VDD VSS n327 NOR2X1 
XU331 n330 n331 VDD VSS n329 NAND2X1 
XU332 N17 n293 VDD VSS n331 NAND2X1 
XU333 N11 VDD VSS n293 INVX1 
XU334 N43 n332 VDD VSS n330 NAND2X1 
XU335 N37 VDD VSS n332 INVX1 
XU336 n333 n334 VDD VSS n328 NAND2X1 
XU337 N108 n335 VDD VSS n334 NAND2X1 
XU338 N102 VDD VSS n335 INVX1 
XU339 n324 n336 VDD VSS n333 NOR2X1 
XU340 N1 n272 VDD VSS n336 NOR2X1 
XU341 N4 VDD VSS n272 INVX1 
XU342 N24 n247 VDD VSS n324 NOR2X1 
XU343 N30 VDD VSS n247 INVX1 
XU344 n337 n338 VDD VSS n326 NOR2X1 
XU345 n339 n340 VDD VSS n338 NAND2X1 
XU346 N82 n341 VDD VSS n340 NAND2X1 
XU347 N76 VDD VSS n341 INVX1 
XU348 N95 n342 VDD VSS n339 NAND2X1 
XU349 N89 VDD VSS n342 INVX1 
XU350 n343 n344 VDD VSS n337 NAND2X1 
XU351 N56 n345 VDD VSS n344 NAND2X1 
XU352 N50 VDD VSS n345 INVX1 
XU353 N69 n346 VDD VSS n343 NAND2X1 
XU354 N63 VDD VSS n346 INVX1 
.ENDS

