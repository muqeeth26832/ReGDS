// SPICE2Verilog Conversion

module c6288 ( N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, N188, N205, N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, N392, N409, N426, N443, N460, N477, N494, N511, N528, N545, N1581, N1901, N2223, N2548, N2877, N3211, N3552, N3895, N4241, N4591, N4946, N5308, N5672, N5971, N6123, N6150, N6160, N6170, N6180, N6190, N6200, N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280, N6287, N6288, VDD, VSS ); 

input N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, N188, N205, N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, N392, N409, N426, N443, N460, N477, N494, N511, N528;
output N545, N1581, N1901, N2223, N2548, N2877, N3211, N3552, N3895, N4241, N4591, N4946, N5308, N5672, N5971, N6123, N6150, N6160, N6170, N6180, N6190, N6200, N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280, N6287, N6288;
inout VDD, VSS;
wire n2209, n2210, n2202, n2242, n2243, n2245, n2267, n2274, n2272, n2248, n2249, n2285, n2283, n2282, n2261, n2260, n2296, n2302, n2304, n2279, n2278, n2322, n2289, n2290, n2331, n2294, n2293, n2301, n2300, n2342, n2348, n2350, n2312, n2311, n2352, n2358, n2360, n2327, n2326, n2378, n2335, n2336, n2389, n2340, n2339, n2347, n2346, n2400, n2406, n2408, n2357, n2356, n2410, n2416, n2418, n2368, n2367, n2420, n2426, n2428, n2383, n2382, n2446, n2393, n2394, n2459, n2398, n2397, n2405, n2404, n2470, n2476, n2478, n2415, n2414, n2480, n2486, n2488, n2425, n2424, n2490, n2496, n2498, n2436, n2435, n2500, n2506, n2508, n2451, n2450, n2526, n2222, n2221, n2203, n2231, n2232, n2230, n2215, n2286, n2284, n2298, n2332, n2330, n2344, n2390, n2388, n2402, n2412, n2422, n2460, n2458, n2474, n2475, n2472, n2484, n2485, n2482, n2494, n2495, n2492, n2204, n2201, n2211, n2212, n2244, n2216, n2220, n2217, n2223, n2224, n2227, n2247, n2246, n2239, n2254, n2252, n2235, n2263, n2255, n2277, n2276, n2307, n2306, n2262, n2280, n2281, n2295, n2258, n2305, n2314, n2325, n2324, n2318, n2363, n2362, n2313, n2353, n2328, n2341, n2292, n2309, n2361, n2370, n2381, n2380, n2374, n2431, n2430, n2369, n2385, n2421, n2384, n2411, n2386, n2399, n2338, n2355, n2419, n2365, n2429, n2438, n2449, n2448, n2442, n2511, n2510, n2437, n2501, n2452, n2491, n2454, n2481, n2456, n2469, n2396, n2433, n2509, n2518, n2529, n2528, n2522, n2205, n2206, n2214, n2228, n2226, n2251, n2259, n2265, n2266, n2264, n2268, n2236, n2275, n2271, n2310, n2316, n2317, n2315, n2319, n2329, n2303, n2366, n2372, n2373, n2371, n2375, n2359, n2387, n2349, n2434, n2440, n2441, n2439, n2443, n2453, n2427, n2455, n2417, n2457, n2407, n2517, n2514, n2520, n2521, n2519, n2523, n2532, n2533, n2507, n2199, n2200, n2207, n2208, n2213, n2219, n2218, n2225, n2229, n2233, n2234, n2237, n2238, n2240, n2241, n2250, n2253, n2256, n2257, n2269, n2270, n2273, n2287, n2288, n2291, n2297, n2299, n2308, n2320, n2321, n2323, n2333, n2334, n2337, n2343, n2345, n2351, n2354, n2364, n2376, n2377, n2379, n2391, n2392, n2395, n2401, n2403, n2409, n2413, n2423, n2432, n2444, n2445, n2447, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2471, n2473, n2477, n2479, n2483, n2487, n2489, n2493, n2497, n2499, n2502, n2503, n2504, n2505, n2512, n2513, n2515, n2516, n2524, n2525, n2527, n2530, n2531, n2541, n2552, n2558, n2560, n2562, n2568, n2570, n2572, n2578, n2580, n2582, n2588, n2590, n2592, n2598, n2600, n2618, n2545, n2546, n2635, n2550, n2549, n2557, n2556, n2646, n2652, n2654, n2567, n2566, n2656, n2662, n2664, n2577, n2576, n2666, n2672, n2674, n2587, n2586, n2676, n2682, n2684, n2597, n2596, n2686, n2692, n2694, n2608, n2607, n2696, n2702, n2704, n2623, n2622, n2722, n2639, n2640, n2741, n2644, n2643, n2651, n2650, n2752, n2758, n2760, n2661, n2660, n2762, n2768, n2770, n2671, n2670, n2772, n2778, n2780, n2681, n2680, n2782, n2788, n2790, n2691, n2690, n2792, n2798, n2800, n2701, n2700, n2802, n2808, n2810, n2712, n2711, n2812, n2818, n2820, n2542, n2540, n2554, n2564, n2574, n2584, n2594, n2636, n2634, n2648, n2658, n2668, n2678, n2688, n2742, n2740, n2756, n2757, n2754, n2766, n2767, n2764, n2776, n2777, n2774, n2786, n2787, n2784, n2796, n2797, n2794, n2806, n2807, n2804, n2816, n2817, n2814, n2593, n2583, n2534, n2573, n2536, n2563, n2538, n2551, n2591, n2601, n2610, n2602, n2621, n2620, n2614, n2707, n2706, n2609, n2697, n2624, n2687, n2626, n2677, n2628, n2667, n2630, n2657, n2632, n2645, n2548, n2605, n2705, n2714, n2725, n2724, n2718, n2823, n2822, n2713, n2729, n2813, n2728, n2803, n2730, n2793, n2732, n2783, n2734, n2773, n2736, n2763, n2738, n2751, n2642, n2699, n2811, n2709, n2821, n2830, n2535, n2537, n2539, n2606, n2612, n2613, n2611, n2615, n2625, n2599, n2627, n2589, n2629, n2579, n2631, n2569, n2633, n2559, n2710, n2716, n2717, n2715, n2719, n2703, n2731, n2693, n2733, n2683, n2735, n2673, n2737, n2663, n2739, n2653, n2829, n2826, n2832, n2833, n2831, n2834, n2835, n2727, n2543, n2544, n2547, n2553, n2555, n2561, n2565, n2571, n2575, n2581, n2585, n2595, n2603, n2604, n2616, n2617, n2619, n2637, n2638, n2641, n2647, n2649, n2655, n2659, n2665, n2669, n2675, n2679, n2685, n2689, n2695, n2698, n2708, n2720, n2721, n2723, n2726, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2753, n2755, n2759, n2761, n2765, n2769, n2771, n2775, n2779, n2781, n2785, n2789, n2791, n2795, n2799, n2801, n2805, n2809, n2815, n2819, n2824, n2825, n2827, n2828, n2836, n2837, n2838, n2859, n2870, n2876, n2878, n2880, n2886, n2888, n2890, n2896, n2898, n2900, n2906, n2908, n2910, n2916, n2918, n2920, n2926, n2928, n2930, n2936, n2938, n2940, n2946, n2948, n2843, n2842, n2966, n2863, n2864, n2989, n2868, n2867, n2875, n2874, n3000, n3006, n3008, n2885, n2884, n3010, n3016, n3018, n2895, n2894, n3020, n3026, n3028, n2905, n2904, n3030, n3036, n3038, n2915, n2914, n3040, n3046, n3048, n2925, n2924, n3050, n3056, n3058, n2935, n2934, n3060, n3066, n3068, n2945, n2944, n3070, n3076, n3078, n2956, n2955, n3080, n3086, n3088, n2971, n2970, n3106, n2993, n2994, n3131, n2860, n2858, n2872, n2882, n2892, n2902, n2912, n2922, n2932, n2990, n2988, n3004, n3005, n3002, n3014, n3015, n3012, n3024, n3025, n3022, n3034, n3035, n3032, n3044, n3045, n3042, n3054, n3055, n3052, n3064, n3065, n3062, n3074, n3075, n3072, n3084, n3085, n3082, n3132, n3130, n2951, n2950, n2941, n2844, n2931, n2846, n2921, n2848, n2911, n2850, n2901, n2852, n2891, n2854, n2881, n2856, n2869, n2949, n2840, n2958, n2969, n2968, n2962, n3091, n3090, n2957, n2973, n3081, n2972, n3071, n2974, n3061, n2976, n3051, n2978, n3041, n2980, n3031, n2982, n3021, n2984, n3011, n2986, n2999, n2866, n2943, n3079, n2953, n3089, n3098, n3109, n3108, n3102, n2845, n2847, n2849, n2851, n2853, n2855, n2857, n2954, n2960, n2961, n2959, n2963, n2947, n2975, n2937, n2977, n2927, n2979, n2917, n2981, n2907, n2983, n2897, n2985, n2887, n2987, n2877, n3097, n3094, n3100, n3101, n3099, n3103, n3112, n3113, n3087, n3114, n3115, n3077, n3116, n3117, n3067, n3118, n3119, n3057, n3120, n3121, n3047, n3122, n3123, n3037, n3124, n3125, n3027, n3126, n3127, n3017, n3128, n3129, n3007, n2839, n2841, n2861, n2862, n2865, n2871, n2873, n2879, n2883, n2889, n2893, n2899, n2903, n2909, n2913, n2919, n2923, n2929, n2933, n2939, n2942, n2952, n2964, n2965, n2967, n2991, n2992, n2995, n2996, n2997, n2998, n3001, n3003, n3009, n3013, n3019, n3023, n3029, n3033, n3039, n3043, n3049, n3053, n3059, n3063, n3069, n3073, n3083, n3092, n3093, n3095, n3096, n3104, n3105, n3107, n3110, n3111, n3133, n3134, n3135, n3136, n3137, n3138, n3142, n3148, n3150, n3152, n3158, n3160, n3162, n3168, n3170, n3172, n3178, n3180, n3182, n3188, n3190, n3192, n3198, n3200, n3202, n3208, n3210, n3212, n3218, n3220, n3222, n3228, n3230, n3232, n3238, n3240, n3258, n3285, n3140, n3139, n3147, n3146, n3292, n3298, n3300, n3157, n3156, n3302, n3308, n3310, n3167, n3166, n3312, n3318, n3320, n3177, n3176, n3322, n3328, n3330, n3187, n3186, n3332, n3338, n3340, n3197, n3196, n3342, n3348, n3350, n3207, n3206, n3352, n3358, n3360, n3217, n3216, n3362, n3368, n3370, n3227, n3226, n3372, n3378, n3380, n3237, n3236, n3382, n3388, n3390, n3248, n3247, n3392, n3398, n3400, n3263, n3262, n3412, n3144, n3154, n3164, n3174, n3184, n3194, n3204, n3214, n3224, n3234, n3286, n3284, n3296, n3297, n3294, n3306, n3307, n3304, n3316, n3317, n3314, n3326, n3327, n3324, n3336, n3337, n3334, n3346, n3347, n3344, n3356, n3357, n3354, n3366, n3367, n3364, n3386, n3387, n3384, n3396, n3397, n3394, n3402, n3403, n3245, n3141, n3241, n3250, n3242, n3261, n3260, n3254, n3393, n3264, n3383, n3266, n3373, n3268, n3363, n3270, n3353, n3272, n3343, n3274, n3333, n3276, n3323, n3278, n3313, n3280, n3303, n3282, n3291, n3401, n3414, n3408, n3415, n3377, n3376, n3424, n3249, n3246, n3252, n3253, n3251, n3255, n3265, n3239, n3267, n3229, n3269, n3219, n3271, n3209, n3273, n3199, n3275, n3189, n3277, n3179, n3279, n3169, n3281, n3159, n3283, n3149, n3406, n3407, n3405, n3409, n3416, n3417, n3419, n3420, n3399, n3421, n3422, n3389, n3423, n3379, n3425, n3426, n3369, n3427, n3428, n3359, n3429, n3430, n3349, n3431, n3432, n3339, n3143, n3145, n3151, n3153, n3155, n3161, n3163, n3165, n3171, n3173, n3175, n3181, n3183, n3185, n3191, n3193, n3195, n3201, n3203, n3205, n3211, n3213, n3215, n3221, n3223, n3225, n3231, n3233, n3235, n3243, n3244, n3256, n3257, n3259, n3287, n3288, n3289, n3290, n3293, n3295, n3299, n3301, n3305, n3309, n3311, n3315, n3319, n3321, n3325, n3329, n3331, n3335, n3341, n3345, n3351, n3355, n3361, n3365, n3371, n3374, n3375, n3381, n3385, n3391, n3395, n3404, n3410, n3411, n3413, n3418, n3445, n3444, n3447, n3455, n3454, n3458, n3464, n3466, n3468, n3474, n3476, n3478, n3484, n3486, n3488, n3494, n3496, n3498, n3504, n3506, n3508, n3514, n3516, n3518, n3524, n3526, n3528, n3534, n3536, n3538, n3544, n3546, n3548, n3554, n3556, n3608, n3607, n3452, n3451, n3610, n3616, n3615, n3463, n3462, n3618, n3626, n3625, n3473, n3472, n3628, n3634, n3636, n3483, n3482, n3638, n3644, n3646, n3493, n3492, n3648, n3654, n3656, n3503, n3502, n3658, n3664, n3666, n3513, n3512, n3668, n3674, n3676, n3523, n3522, n3678, n3684, n3686, n3533, n3532, n3688, n3694, n3696, n3543, n3542, n3698, n3704, n3706, n3553, n3552, n3708, n3714, n3716, n3449, n3460, n3470, n3480, n3490, n3500, n3510, n3520, n3540, n3550, n3560, n3561, n3559, n3622, n3623, n3620, n3632, n3633, n3630, n3642, n3643, n3640, n3652, n3653, n3650, n3662, n3663, n3660, n3672, n3673, n3670, n3682, n3683, n3680, n3692, n3693, n3690, n3702, n3703, n3700, n3720, n3721, n3719, n3499, n3489, n3433, n3479, n3435, n3469, n3437, n3459, n3439, n3443, n3441, n3446, n3457, n3537, n3562, n3558, n3570, n3569, n3568, n3578, n3579, n3726, n3725, n3718, n3581, n3709, n3583, n3586, n3699, n3585, n3689, n3587, n3679, n3589, n3669, n3591, n3659, n3593, n3649, n3595, n3639, n3597, n3629, n3599, n3619, n3601, n3604, n3605, n3609, n3606, n3450, n3617, n3461, n3627, n3531, n3697, n3580, n3722, n3434, n3436, n3438, n3440, n3442, n3456, n3565, n3567, n3577, n3575, n3563, n3582, n3555, n3584, n3545, n3535, n3588, n3525, n3590, n3515, n3592, n3505, n3594, n3495, n3596, n3485, n3598, n3475, n3600, n3465, n3602, n3453, n3603, n3448, n3467, n3471, n3477, n3481, n3487, n3491, n3497, n3501, n3507, n3509, n3511, n3517, n3519, n3521, n3527, n3529, n3530, n3539, n3541, n3547, n3549, n3551, n3557, n3564, n3566, n3571, n3572, n3573, n3574, n3576, n3611, n3612, n3613, n3614, n3621, n3624, n3631, n3635, n3637, n3641, n3645, n3647, n3651, n3655, n3657, n3661, n3665, n3667, n3671, n3675, n3677, n3681, n3685, n3687, n3691, n3695, n3701, n3705, n3707, n3710, n3711, n3712, n3713, n3715, n3717, n3723, n3724, n3727, n3775, n3783, n3782, n3785, n3793, n3792, n3795, n3801, n3803, n3805, n3811, n3813, n3815, n3821, n3823, n3825, n3831, n3833, n3835, n3841, n3843, n3845, n3851, n3853, n3855, n3861, n3863, n3865, n3871, n3873, n3928, n3780, n3790, n3789, n3931, n3925, n3938, n3800, n3799, n3940, n3921, n3947, n3810, n3809, n3949, n3955, n3957, n3820, n3819, n3959, n3965, n3967, n3830, n3829, n3969, n3975, n3977, n3840, n3839, n3979, n3985, n3987, n3850, n3849, n3989, n3995, n3997, n3860, n3859, n3999, n4005, n4007, n3870, n3869, n4009, n4015, n4017, n3779, n3777, n3857, n3877, n3878, n3876, n3893, n3736, n3892, n3935, n3936, n3933, n4003, n4004, n4001, n4021, n4022, n4020, n3730, n3729, n3728, n3735, n3733, n3737, n3747, n3748, n3883, n3882, n3751, n3875, n3750, n3866, n3752, n3856, n3754, n3846, n3756, n3836, n3758, n3826, n3760, n3816, n3762, n3806, n3764, n3796, n3766, n3786, n3768, n3774, n3772, n3784, n3794, n3874, n3749, n3879, n3887, n3886, n3885, n3890, n3897, n3901, n3902, n4027, n4026, n3905, n4019, n3904, n4010, n3906, n3909, n4000, n3908, n3911, n3990, n3910, n3913, n3980, n3912, n3915, n3970, n3914, n3917, n3960, n3916, n3920, n3950, n3918, n3924, n3941, n3922, n3932, n3926, n3778, n3930, n3788, n3939, n3798, n3948, n3808, n3958, n3818, n3968, n3828, n3978, n3838, n3988, n3848, n3998, n3868, n4018, n3903, n4023, n3732, n3740, n3742, n3738, n3743, n3744, n3745, n3746, n3753, n3755, n3757, n3759, n3761, n3763, n3765, n3767, n3769, n3771, n3884, n3889, n3898, n3880, n3872, n3907, n3862, n3852, n3842, n3832, n3822, n3812, n3919, n3802, n3923, n3791, n3927, n3781, n3929, n3731, n3734, n3739, n3741, n3770, n3773, n3776, n3787, n3797, n3804, n3807, n3814, n3817, n3824, n3827, n3834, n3837, n3844, n3847, n3854, n3858, n3864, n3867, n3881, n3888, n3891, n3895, n3896, n3894, n3899, n3900, n3934, n3937, n3942, n3943, n3944, n3945, n3946, n3951, n3952, n3953, n3954, n3956, n3961, n3962, n3963, n3964, n3966, n3971, n3972, n3973, n3974, n3976, n3981, n3982, n3983, n3984, n3986, n3991, n3992, n3993, n3994, n3996, n4002, n4006, n4008, n4011, n4012, n4013, n4014, n4016, n4024, n4025, n4028, n4069, n4071, n4066, n4078, n4080, n4062, n4087, n4089, n4095, n4097, n4099, n4105, n4107, n4109, n4115, n4117, n4119, n4125, n4127, n4129, n4135, n4137, n4139, n4145, n4147, n4196, n4076, n4085, n4084, n4198, n4193, n4205, n4094, n4093, n4207, n4189, n4214, n4104, n4103, n4216, n4222, n4224, n4114, n4113, n4226, n4232, n4234, n4124, n4123, n4236, n4242, n4244, n4134, n4133, n4246, n4252, n4254, n4144, n4143, n4256, n4262, n4264, n4312, n4203, n4212, n4211, n4314, n4309, n4321, n4075, n4073, n4131, n4151, n4152, n4150, n4167, n4037, n4166, n4202, n4200, n4250, n4251, n4248, n4268, n4269, n4267, n4318, n4319, n4316, n4031, n4030, n4029, n4036, n4034, n4041, n4044, n4045, n4157, n4156, n4048, n4149, n4047, n4140, n4049, n4052, n4130, n4051, n4054, n4120, n4053, n4056, n4110, n4055, n4058, n4100, n4057, n4061, n4090, n4059, n4065, n4081, n4063, n4072, n4067, n4070, n4079, n4088, n4098, n4108, n4118, n4128, n4148, n4046, n4153, n4161, n4160, n4159, n4164, n4170, n4173, n4174, n4274, n4273, n4177, n4266, n4176, n4257, n4178, n4181, n4247, n4180, n4183, n4237, n4182, n4185, n4227, n4184, n4188, n4217, n4186, n4192, n4208, n4190, n4199, n4194, n4074, n4197, n4083, n4206, n4092, n4215, n4102, n4225, n4112, n4235, n4122, n4245, n4142, n4265, n4175, n4270, n4278, n4277, n4276, n4283, n4281, n4288, n4291, n4292, n4261, n4260, n4295, n4241, n4240, n4299, n4231, n4230, n4301, n4308, n4315, n4310, n4201, n4313, n4033, n4050, n4060, n4064, n4068, n4158, n4163, n4154, n4146, n4179, n4136, n4126, n4116, n4106, n4187, n4096, n4191, n4086, n4195, n4077, n4275, n4280, n4271, n4294, n4263, n4296, n4297, n4253, n4298, n4243, n4300, n4233, n4302, n4303, n4223, n4304, n4305, n4306, n4307, n4213, n4311, n4204, n4032, n4035, n4038, n4039, n4040, n4042, n4043, n4082, n4091, n4101, n4111, n4121, n4132, n4138, n4141, n4155, n4162, n4165, n4168, n4169, n4171, n4172, n4209, n4210, n4218, n4219, n4220, n4221, n4228, n4229, n4238, n4239, n4249, n4255, n4258, n4259, n4272, n4279, n4282, n4284, n4285, n4286, n4287, n4289, n4290, n4317, n4320, n4293, n4323, n4330, n4332, n4338, n4340, n4342, n4348, n4350, n4352, n4358, n4360, n4362, n4368, n4370, n4415, n4328, n4327, n4417, n4412, n4424, n4337, n4336, n4426, n4408, n4433, n4347, n4346, n4435, n4441, n4443, n4357, n4356, n4445, n4451, n4453, n4367, n4366, n4455, n4461, n4463, n4507, n4422, n4431, n4430, n4509, n4504, n4516, n4440, n4439, n4518, n4500, n4525, n4450, n4449, n4527, n4533, n4535, n4460, n4459, n4537, n4543, n4545, n4584, n4514, n4523, n4522, n4586, n4581, n4593, n4532, n4531, n4595, n4603, n4602, n4542, n4541, n4605, n4611, n4613, n4354, n4374, n4375, n4373, n4390, n4389, n4421, n4419, n4447, n4467, n4468, n4466, n4513, n4511, n4529, n4549, n4550, n4548, n4565, n4483, n4564, n4590, n4591, n4588, n4599, n4600, n4597, n4331, n4341, n4351, n4371, n4376, n4372, n4384, n4383, n4382, n4387, n4393, n4396, n4397, n4473, n4472, n4400, n4465, n4399, n4456, n4401, n4404, n4446, n4403, n4407, n4436, n4405, n4411, n4427, n4409, n4418, n4413, n4416, n4326, n4425, n4335, n4434, n4345, n4444, n4365, n4464, n4398, n4469, n4477, n4476, n4475, n4482, n4480, n4487, n4490, n4491, n4555, n4554, n4494, n4547, n4493, n4538, n4495, n4499, n4528, n4497, n4503, n4519, n4501, n4510, n4505, n4420, n4508, n4429, n4517, n4438, n4526, n4458, n4546, n4492, n4551, n4559, n4558, n4557, n4562, n4568, n4571, n4572, n4575, n4616, n4615, n4574, n4606, n4576, n4580, n4596, n4578, n4587, n4582, n4512, n4585, n4521, n4594, n4530, n4604, n4540, n4614, n4379, n4381, n4386, n4377, n4369, n4402, n4359, n4349, n4406, n4339, n4410, n4329, n4414, n4474, n4479, n4470, n4462, n4496, n4452, n4498, n4442, n4502, n4432, n4506, n4423, n4556, n4561, n4552, n4544, n4577, n4534, n4579, n4524, n4583, n4515, n4322, n4324, n4325, n4333, n4334, n4343, n4344, n4353, n4355, n4361, n4363, n4364, n4378, n4380, n4385, n4388, n4391, n4392, n4394, n4395, n4428, n4437, n4448, n4454, n4457, n4471, n4478, n4481, n4484, n4485, n4486, n4488, n4489, n4520, n4536, n4539, n4553, n4560, n4563, n4566, n4567, n4569, n4570, n4589, n4592, n4598, n4601, n4607, n4608, n4609, n4610, n4612, n4573, n4651, n4653, n4661, n4660, n4663, n4646, n4670, n4705, n4658, n4668, n4667, n4707, n4702, n4714, n4746, n4712, n4657, n4655, n4674, n4675, n4673, n4690, n4633, n4689, n4711, n4709, n4718, n4719, n4717, n4766, n4734, n4765, n4780, n4779, n4751, n4619, n4627, n4626, n4625, n4632, n4630, n4637, n4640, n4641, n4680, n4679, n4617, n4645, n4672, n4643, n4664, n4647, n4654, n4649, n4652, n4662, n4671, n4642, n4676, n4684, n4683, n4682, n4687, n4693, n4696, n4697, n4724, n4723, n4701, n4716, n4699, n4708, n4703, n4656, n4706, n4666, n4715, n4698, n4720, n4728, n4727, n4726, n4733, n4731, n4738, n4741, n4742, n4756, n4755, n4749, n4748, n4744, n4710, n4747, n4743, n4752, n4760, n4759, n4758, n4763, n4769, n4772, n4773, n4750, n4753, n4778, n4776, n4781, n4782, n4787, n4785, n4792, n4788, n4799, n4797, n4808, n4809, n4800, n4622, n4624, n4629, n4618, n4620, n4644, n4648, n4650, n4681, n4686, n4677, n4700, n4669, n4704, n4659, n4725, n4730, n4721, n4745, n4713, n4757, n4762, n4775, n4784, n4796, n4806, n4807, n4621, n4623, n4628, n4631, n4634, n4635, n4636, n4638, n4639, n4665, n4678, n4685, n4688, n4691, n4692, n4694, n4695, n4722, n4729, n4732, n4735, n4736, n4737, n4739, n4740, n4754, n4761, n4764, n4767, n4768, n4770, n4771, n4774, n4777, n4783, n4786, n4789, n4790, n4791, n4793, n4794, n4795, n4798, n4801, n4802, n4803, n4804, n4805;

XOR2 X1 (.A(n2209), .B(n2210), .Y(n2202), .VDD(VDD), .GND(VSS) );
XOR2 X2 (.A(n2242), .B(n2243), .Y(n2245), .VDD(VDD), .GND(VSS) );
XOR2 X3 (.A(n2267), .B(n2274), .Y(n2272), .VDD(VDD), .GND(VSS) );
XOR2 X4 (.A(n2248), .B(n2249), .Y(n2285), .VDD(VDD), .GND(VSS) );
XOR2 X5 (.A(n2283), .B(n2282), .Y(n2248), .VDD(VDD), .GND(VSS) );
XOR2 X6 (.A(n2261), .B(n2260), .Y(n2296), .VDD(VDD), .GND(VSS) );
XOR2 X7 (.A(n2302), .B(n2261), .Y(n2304), .VDD(VDD), .GND(VSS) );
XOR2 X8 (.A(n2279), .B(n2278), .Y(n2322), .VDD(VDD), .GND(VSS) );
XOR2 X9 (.A(n2289), .B(n2290), .Y(n2331), .VDD(VDD), .GND(VSS) );
XOR2 X10 (.A(n2294), .B(n2293), .Y(n2289), .VDD(VDD), .GND(VSS) );
XOR2 X11 (.A(n2301), .B(n2300), .Y(n2342), .VDD(VDD), .GND(VSS) );
XOR2 X12 (.A(n2300), .B(n2348), .Y(n2350), .VDD(VDD), .GND(VSS) );
XOR2 X13 (.A(n2312), .B(n2311), .Y(n2352), .VDD(VDD), .GND(VSS) );
XOR2 X14 (.A(n2358), .B(n2312), .Y(n2360), .VDD(VDD), .GND(VSS) );
XOR2 X15 (.A(n2327), .B(n2326), .Y(n2378), .VDD(VDD), .GND(VSS) );
XOR2 X16 (.A(n2335), .B(n2336), .Y(n2389), .VDD(VDD), .GND(VSS) );
XOR2 X17 (.A(n2340), .B(n2339), .Y(n2335), .VDD(VDD), .GND(VSS) );
XOR2 X18 (.A(n2347), .B(n2346), .Y(n2400), .VDD(VDD), .GND(VSS) );
XOR2 X19 (.A(n2346), .B(n2406), .Y(n2408), .VDD(VDD), .GND(VSS) );
XOR2 X20 (.A(n2357), .B(n2356), .Y(n2410), .VDD(VDD), .GND(VSS) );
XOR2 X21 (.A(n2416), .B(n2357), .Y(n2418), .VDD(VDD), .GND(VSS) );
XOR2 X22 (.A(n2368), .B(n2367), .Y(n2420), .VDD(VDD), .GND(VSS) );
XOR2 X23 (.A(n2426), .B(n2368), .Y(n2428), .VDD(VDD), .GND(VSS) );
XOR2 X24 (.A(n2383), .B(n2382), .Y(n2446), .VDD(VDD), .GND(VSS) );
XOR2 X25 (.A(n2393), .B(n2394), .Y(n2459), .VDD(VDD), .GND(VSS) );
XOR2 X26 (.A(n2398), .B(n2397), .Y(n2393), .VDD(VDD), .GND(VSS) );
XOR2 X27 (.A(n2405), .B(n2404), .Y(n2470), .VDD(VDD), .GND(VSS) );
XOR2 X28 (.A(n2404), .B(n2476), .Y(n2478), .VDD(VDD), .GND(VSS) );
XOR2 X29 (.A(n2415), .B(n2414), .Y(n2480), .VDD(VDD), .GND(VSS) );
XOR2 X30 (.A(n2414), .B(n2486), .Y(n2488), .VDD(VDD), .GND(VSS) );
XOR2 X31 (.A(n2425), .B(n2424), .Y(n2490), .VDD(VDD), .GND(VSS) );
XOR2 X32 (.A(n2424), .B(n2496), .Y(n2498), .VDD(VDD), .GND(VSS) );
XOR2 X33 (.A(n2436), .B(n2435), .Y(n2500), .VDD(VDD), .GND(VSS) );
XOR2 X34 (.A(n2506), .B(n2436), .Y(n2508), .VDD(VDD), .GND(VSS) );
XOR2 X35 (.A(n2451), .B(n2450), .Y(n2526), .VDD(VDD), .GND(VSS) );
OR2X1 X36 (.A(n2222), .B(n2221), .VDD(VDD), .VSS(VSS), .Y(n2203) );
OR2X1 X37 (.A(n2231), .B(n2232), .VDD(VDD), .VSS(VSS), .Y(n2230) );
OR2X1 X38 (.A(n2243), .B(n2242), .VDD(VDD), .VSS(VSS), .Y(n2215) );
OR2X1 X39 (.A(n2285), .B(n2286), .VDD(VDD), .VSS(VSS), .Y(n2284) );
OR2X1 X40 (.A(n2300), .B(n2301), .VDD(VDD), .VSS(VSS), .Y(n2298) );
OR2X1 X41 (.A(n2331), .B(n2332), .VDD(VDD), .VSS(VSS), .Y(n2330) );
OR2X1 X42 (.A(n2346), .B(n2347), .VDD(VDD), .VSS(VSS), .Y(n2344) );
OR2X1 X43 (.A(n2389), .B(n2390), .VDD(VDD), .VSS(VSS), .Y(n2388) );
OR2X1 X44 (.A(n2404), .B(n2405), .VDD(VDD), .VSS(VSS), .Y(n2402) );
OR2X1 X45 (.A(n2414), .B(n2415), .VDD(VDD), .VSS(VSS), .Y(n2412) );
OR2X1 X46 (.A(n2424), .B(n2425), .VDD(VDD), .VSS(VSS), .Y(n2422) );
OR2X1 X47 (.A(n2459), .B(n2460), .VDD(VDD), .VSS(VSS), .Y(n2458) );
OR2X1 X48 (.A(n2474), .B(n2475), .VDD(VDD), .VSS(VSS), .Y(n2472) );
OR2X1 X49 (.A(n2484), .B(n2485), .VDD(VDD), .VSS(VSS), .Y(n2482) );
OR2X1 X50 (.A(n2494), .B(n2495), .VDD(VDD), .VSS(VSS), .Y(n2492) );
AND2X1 X51 (.A(n2203), .B(n2204), .VDD(VDD), .VSS(VSS), .Y(n2201) );
AND2X1 X52 (.A(n2211), .B(n2212), .VDD(VDD), .VSS(VSS), .Y(n2210) );
AND2X1 X53 (.A(n2244), .B(n2245), .VDD(VDD), .VSS(VSS), .Y(n2216) );
AND2X1 X54 (.A(n2203), .B(n2220), .VDD(VDD), .VSS(VSS), .Y(n2217) );
AND2X1 X55 (.A(n2223), .B(n2224), .VDD(VDD), .VSS(VSS), .Y(n2221) );
AND2X1 X56 (.A(n2211), .B(n2230), .VDD(VDD), .VSS(VSS), .Y(n2227) );
AND2X1 X57 (.A(n2247), .B(n2246), .VDD(VDD), .VSS(VSS), .Y(n2239) );
AND2X1 X58 (.A(n2254), .B(n2223), .VDD(VDD), .VSS(VSS), .Y(n2252) );
AND2X1 X59 (.A(n2235), .B(n2263), .VDD(VDD), .VSS(VSS), .Y(n2255) );
AND2X1 X60 (.A(n2277), .B(n2276), .VDD(VDD), .VSS(VSS), .Y(n2267) );
AND2X1 X61 (.A(n2307), .B(n2306), .VDD(VDD), .VSS(VSS), .Y(n2262) );
AND2X1 X62 (.A(n2280), .B(n2281), .VDD(VDD), .VSS(VSS), .Y(n2242) );
AND2X1 X63 (.A(n2295), .B(n2281), .VDD(VDD), .VSS(VSS), .Y(n2282) );
AND2X1 X64 (.A(n2258), .B(n2305), .VDD(VDD), .VSS(VSS), .Y(n2260) );
AND2X1 X65 (.A(n2276), .B(n2314), .VDD(VDD), .VSS(VSS), .Y(n2306) );
AND2X1 X66 (.A(n2325), .B(n2324), .VDD(VDD), .VSS(VSS), .Y(n2318) );
AND2X1 X67 (.A(n2363), .B(n2362), .VDD(VDD), .VSS(VSS), .Y(n2313) );
AND2X1 X68 (.A(n2353), .B(n2352), .VDD(VDD), .VSS(VSS), .Y(n2328) );
AND2X1 X69 (.A(n2341), .B(n2292), .VDD(VDD), .VSS(VSS), .Y(n2293) );
AND2X1 X70 (.A(N511), .B(N205), .VDD(VDD), .VSS(VSS), .Y(n2301) );
AND2X1 X71 (.A(n2309), .B(n2361), .VDD(VDD), .VSS(VSS), .Y(n2311) );
AND2X1 X72 (.A(n2324), .B(n2370), .VDD(VDD), .VSS(VSS), .Y(n2362) );
AND2X1 X73 (.A(n2381), .B(n2380), .VDD(VDD), .VSS(VSS), .Y(n2374) );
AND2X1 X74 (.A(n2431), .B(n2430), .VDD(VDD), .VSS(VSS), .Y(n2369) );
AND2X1 X75 (.A(n2357), .B(n2356), .VDD(VDD), .VSS(VSS), .Y(n2385) );
AND2X1 X76 (.A(n2421), .B(n2420), .VDD(VDD), .VSS(VSS), .Y(n2384) );
AND2X1 X77 (.A(n2411), .B(n2410), .VDD(VDD), .VSS(VSS), .Y(n2386) );
AND2X1 X78 (.A(n2399), .B(n2338), .VDD(VDD), .VSS(VSS), .Y(n2339) );
AND2X1 X79 (.A(N511), .B(N188), .VDD(VDD), .VSS(VSS), .Y(n2347) );
AND2X1 X80 (.A(n2355), .B(n2419), .VDD(VDD), .VSS(VSS), .Y(n2356) );
AND2X1 X81 (.A(n2365), .B(n2429), .VDD(VDD), .VSS(VSS), .Y(n2367) );
AND2X1 X82 (.A(n2380), .B(n2438), .VDD(VDD), .VSS(VSS), .Y(n2430) );
AND2X1 X83 (.A(n2449), .B(n2448), .VDD(VDD), .VSS(VSS), .Y(n2442) );
AND2X1 X84 (.A(n2511), .B(n2510), .VDD(VDD), .VSS(VSS), .Y(n2437) );
AND2X1 X85 (.A(n2501), .B(n2500), .VDD(VDD), .VSS(VSS), .Y(n2452) );
AND2X1 X86 (.A(n2491), .B(n2490), .VDD(VDD), .VSS(VSS), .Y(n2454) );
AND2X1 X87 (.A(n2481), .B(n2480), .VDD(VDD), .VSS(VSS), .Y(n2456) );
AND2X1 X88 (.A(n2469), .B(n2396), .VDD(VDD), .VSS(VSS), .Y(n2397) );
AND2X1 X89 (.A(N511), .B(N171), .VDD(VDD), .VSS(VSS), .Y(n2405) );
AND2X1 X90 (.A(N494), .B(N188), .VDD(VDD), .VSS(VSS), .Y(n2415) );
AND2X1 X91 (.A(N477), .B(N205), .VDD(VDD), .VSS(VSS), .Y(n2425) );
AND2X1 X92 (.A(n2433), .B(n2509), .VDD(VDD), .VSS(VSS), .Y(n2435) );
AND2X1 X93 (.A(n2448), .B(n2518), .VDD(VDD), .VSS(VSS), .Y(n2510) );
AND2X1 X94 (.A(n2529), .B(n2528), .VDD(VDD), .VSS(VSS), .Y(n2522) );
NOR2X1 X95 (.A(n2205), .B(n2206), .Y(N6287), .VDD(VDD), .GND(VSS) );
NOR2X1 X96 (.A(n2216), .B(n2217), .Y(n2214), .VDD(VDD), .GND(VSS) );
NOR2X1 X97 (.A(n2227), .B(n2228), .Y(n2226), .VDD(VDD), .GND(VSS) );
NOR2X1 X98 (.A(n2252), .B(n2205), .Y(n2251), .VDD(VDD), .GND(VSS) );
NOR2X1 X99 (.A(n2262), .B(n2255), .Y(n2259), .VDD(VDD), .GND(VSS) );
NOR2X1 X100 (.A(n2265), .B(n2266), .Y(n2264), .VDD(VDD), .GND(VSS) );
NOR2X1 X101 (.A(n2267), .B(n2268), .Y(n2266), .VDD(VDD), .GND(VSS) );
NOR2X1 X102 (.A(N494), .B(n2236), .Y(n2265), .VDD(VDD), .GND(VSS) );
NOR2X1 X103 (.A(n2275), .B(n2271), .Y(n2274), .VDD(VDD), .GND(VSS) );
NOR2X1 X104 (.A(n2313), .B(n2306), .Y(n2310), .VDD(VDD), .GND(VSS) );
NOR2X1 X105 (.A(n2316), .B(n2317), .Y(n2315), .VDD(VDD), .GND(VSS) );
NOR2X1 X106 (.A(n2318), .B(n2319), .Y(n2317), .VDD(VDD), .GND(VSS) );
NOR2X1 X107 (.A(N477), .B(n2279), .Y(n2316), .VDD(VDD), .GND(VSS) );
NOR2X1 X108 (.A(n2328), .B(n2329), .Y(n2303), .VDD(VDD), .GND(VSS) );
NOR2X1 X109 (.A(n2301), .B(n2300), .Y(n2329), .VDD(VDD), .GND(VSS) );
NOR2X1 X110 (.A(n2369), .B(n2362), .Y(n2366), .VDD(VDD), .GND(VSS) );
NOR2X1 X111 (.A(n2372), .B(n2373), .Y(n2371), .VDD(VDD), .GND(VSS) );
NOR2X1 X112 (.A(n2374), .B(n2375), .Y(n2373), .VDD(VDD), .GND(VSS) );
NOR2X1 X113 (.A(N460), .B(n2327), .Y(n2372), .VDD(VDD), .GND(VSS) );
NOR2X1 X114 (.A(n2384), .B(n2385), .Y(n2359), .VDD(VDD), .GND(VSS) );
NOR2X1 X115 (.A(n2386), .B(n2387), .Y(n2349), .VDD(VDD), .GND(VSS) );
NOR2X1 X116 (.A(n2347), .B(n2346), .Y(n2387), .VDD(VDD), .GND(VSS) );
NOR2X1 X117 (.A(n2437), .B(n2430), .Y(n2434), .VDD(VDD), .GND(VSS) );
NOR2X1 X118 (.A(n2440), .B(n2441), .Y(n2439), .VDD(VDD), .GND(VSS) );
NOR2X1 X119 (.A(n2442), .B(n2443), .Y(n2441), .VDD(VDD), .GND(VSS) );
NOR2X1 X120 (.A(N443), .B(n2383), .Y(n2440), .VDD(VDD), .GND(VSS) );
NOR2X1 X121 (.A(n2452), .B(n2453), .Y(n2427), .VDD(VDD), .GND(VSS) );
NOR2X1 X122 (.A(n2425), .B(n2424), .Y(n2453), .VDD(VDD), .GND(VSS) );
NOR2X1 X123 (.A(n2454), .B(n2455), .Y(n2417), .VDD(VDD), .GND(VSS) );
NOR2X1 X124 (.A(n2415), .B(n2414), .Y(n2455), .VDD(VDD), .GND(VSS) );
NOR2X1 X125 (.A(n2456), .B(n2457), .Y(n2407), .VDD(VDD), .GND(VSS) );
NOR2X1 X126 (.A(n2405), .B(n2404), .Y(n2457), .VDD(VDD), .GND(VSS) );
NOR2X1 X127 (.A(n2517), .B(n2510), .Y(n2514), .VDD(VDD), .GND(VSS) );
NOR2X1 X128 (.A(n2520), .B(n2521), .Y(n2519), .VDD(VDD), .GND(VSS) );
NOR2X1 X129 (.A(n2522), .B(n2523), .Y(n2521), .VDD(VDD), .GND(VSS) );
NOR2X1 X130 (.A(N426), .B(n2451), .Y(n2520), .VDD(VDD), .GND(VSS) );
NOR2X1 X131 (.A(n2532), .B(n2533), .Y(n2507), .VDD(VDD), .GND(VSS) );
NAND2X1 X132 (.A(n2199), .B(n2200), .Y(N6288), .VDD(VDD), .GND(VSS) );
NAND2X1 X133 (.A(n2201), .B(n2202), .Y(n2200), .VDD(VDD), .GND(VSS) );
NAND2X1 X134 (.A(N256), .B(n2199), .Y(n2206), .VDD(VDD), .GND(VSS) );
NAND2X1 X135 (.A(n2207), .B(n2208), .Y(n2199), .VDD(VDD), .GND(VSS) );
NAND2X1 X136 (.A(n2204), .B(n2203), .Y(n2208), .VDD(VDD), .GND(VSS) );
NAND2X1 X137 (.A(N528), .B(N256), .Y(n2209), .VDD(VDD), .GND(VSS) );
NAND2X1 X138 (.A(n2204), .B(n2213), .Y(N6280), .VDD(VDD), .GND(VSS) );
NAND2X1 X139 (.A(n2214), .B(n2215), .Y(n2213), .VDD(VDD), .GND(VSS) );
NAND2X1 X140 (.A(n2217), .B(n2219), .Y(n2204), .VDD(VDD), .GND(VSS) );
NAND2X1 X141 (.A(n2215), .B(n2218), .Y(n2219), .VDD(VDD), .GND(VSS) );
NAND2X1 X142 (.A(n2221), .B(n2222), .Y(n2220), .VDD(VDD), .GND(VSS) );
NAND2X1 X143 (.A(n2212), .B(n2225), .Y(n2222), .VDD(VDD), .GND(VSS) );
NAND2X1 X144 (.A(n2226), .B(N528), .Y(n2225), .VDD(VDD), .GND(VSS) );
NAND2X1 X145 (.A(n2227), .B(n2229), .Y(n2212), .VDD(VDD), .GND(VSS) );
NAND2X1 X146 (.A(N528), .B(N239), .Y(n2229), .VDD(VDD), .GND(VSS) );
NAND2X1 X147 (.A(n2231), .B(n2233), .Y(n2211), .VDD(VDD), .GND(VSS) );
NAND2X1 X148 (.A(N256), .B(N511), .Y(n2233), .VDD(VDD), .GND(VSS) );
NAND2X1 X149 (.A(n2234), .B(n2235), .Y(n2231), .VDD(VDD), .GND(VSS) );
NAND2X1 X150 (.A(n2236), .B(n2237), .Y(n2234), .VDD(VDD), .GND(VSS) );
NAND2X1 X151 (.A(N494), .B(N256), .Y(n2237), .VDD(VDD), .GND(VSS) );
NAND2X1 X152 (.A(n2218), .B(n2238), .Y(N6270), .VDD(VDD), .GND(VSS) );
NAND2X1 X153 (.A(n2239), .B(n2240), .Y(n2238), .VDD(VDD), .GND(VSS) );
NAND2X1 X154 (.A(n2215), .B(n2241), .Y(n2240), .VDD(VDD), .GND(VSS) );
NAND2X1 X155 (.A(n2242), .B(n2243), .Y(n2241), .VDD(VDD), .GND(VSS) );
NAND2X1 X156 (.A(n2248), .B(n2249), .Y(n2246), .VDD(VDD), .GND(VSS) );
NAND2X1 X157 (.A(n2224), .B(n2250), .Y(n2243), .VDD(VDD), .GND(VSS) );
NAND2X1 X158 (.A(n2251), .B(N222), .Y(n2250), .VDD(VDD), .GND(VSS) );
NAND2X1 X159 (.A(n2252), .B(n2253), .Y(n2224), .VDD(VDD), .GND(VSS) );
NAND2X1 X160 (.A(N222), .B(N528), .Y(n2253), .VDD(VDD), .GND(VSS) );
NAND2X1 X161 (.A(n2255), .B(n2256), .Y(n2223), .VDD(VDD), .GND(VSS) );
NAND2X1 X162 (.A(n2257), .B(n2258), .Y(n2256), .VDD(VDD), .GND(VSS) );
NAND2X1 X163 (.A(n2259), .B(n2257), .Y(n2254), .VDD(VDD), .GND(VSS) );
NAND2X1 X164 (.A(n2260), .B(n2261), .Y(n2257), .VDD(VDD), .GND(VSS) );
NAND2X1 X165 (.A(n2264), .B(N511), .Y(n2263), .VDD(VDD), .GND(VSS) );
NAND2X1 X166 (.A(n2269), .B(n2270), .Y(n2268), .VDD(VDD), .GND(VSS) );
NAND2X1 X167 (.A(N239), .B(n2271), .Y(n2269), .VDD(VDD), .GND(VSS) );
NAND2X1 X168 (.A(n2272), .B(n2273), .Y(n2235), .VDD(VDD), .GND(VSS) );
NAND2X1 X169 (.A(N511), .B(N239), .Y(n2273), .VDD(VDD), .GND(VSS) );
NAND2X1 X170 (.A(n2278), .B(n2279), .Y(n2277), .VDD(VDD), .GND(VSS) );
NAND2X1 X171 (.A(n2282), .B(n2283), .Y(n2280), .VDD(VDD), .GND(VSS) );
NAND2X1 X172 (.A(n2247), .B(n2284), .Y(N6260), .VDD(VDD), .GND(VSS) );
NAND2X1 X173 (.A(n2285), .B(n2286), .Y(n2247), .VDD(VDD), .GND(VSS) );
NAND2X1 X174 (.A(n2287), .B(n2288), .Y(n2286), .VDD(VDD), .GND(VSS) );
NAND2X1 X175 (.A(n2289), .B(n2290), .Y(n2287), .VDD(VDD), .GND(VSS) );
NAND2X1 X176 (.A(n2291), .B(n2292), .Y(n2249), .VDD(VDD), .GND(VSS) );
NAND2X1 X177 (.A(n2293), .B(n2294), .Y(n2291), .VDD(VDD), .GND(VSS) );
NAND2X1 X178 (.A(n2296), .B(n2297), .Y(n2281), .VDD(VDD), .GND(VSS) );
NAND2X1 X179 (.A(n2298), .B(n2299), .Y(n2297), .VDD(VDD), .GND(VSS) );
NAND2X1 X180 (.A(n2303), .B(n2304), .Y(n2295), .VDD(VDD), .GND(VSS) );
NAND2X1 X181 (.A(N222), .B(N511), .Y(n2261), .VDD(VDD), .GND(VSS) );
NAND2X1 X182 (.A(n2308), .B(n2309), .Y(n2307), .VDD(VDD), .GND(VSS) );
NAND2X1 X183 (.A(n2310), .B(n2308), .Y(n2305), .VDD(VDD), .GND(VSS) );
NAND2X1 X184 (.A(n2311), .B(n2312), .Y(n2308), .VDD(VDD), .GND(VSS) );
NAND2X1 X185 (.A(n2315), .B(N494), .Y(n2314), .VDD(VDD), .GND(VSS) );
NAND2X1 X186 (.A(n2320), .B(n2270), .Y(n2319), .VDD(VDD), .GND(VSS) );
NAND2X1 X187 (.A(N239), .B(n2321), .Y(n2320), .VDD(VDD), .GND(VSS) );
NAND2X1 X188 (.A(n2322), .B(n2323), .Y(n2276), .VDD(VDD), .GND(VSS) );
NAND2X1 X189 (.A(N494), .B(N239), .Y(n2323), .VDD(VDD), .GND(VSS) );
NAND2X1 X190 (.A(N477), .B(N256), .Y(n2278), .VDD(VDD), .GND(VSS) );
NAND2X1 X191 (.A(n2326), .B(n2327), .Y(n2325), .VDD(VDD), .GND(VSS) );
NAND2X1 X192 (.A(N205), .B(N528), .Y(n2283), .VDD(VDD), .GND(VSS) );
NAND2X1 X193 (.A(n2288), .B(n2330), .Y(N6250), .VDD(VDD), .GND(VSS) );
NAND2X1 X194 (.A(n2331), .B(n2332), .Y(n2288), .VDD(VDD), .GND(VSS) );
NAND2X1 X195 (.A(n2333), .B(n2334), .Y(n2332), .VDD(VDD), .GND(VSS) );
NAND2X1 X196 (.A(n2335), .B(n2336), .Y(n2333), .VDD(VDD), .GND(VSS) );
NAND2X1 X197 (.A(n2337), .B(n2338), .Y(n2290), .VDD(VDD), .GND(VSS) );
NAND2X1 X198 (.A(n2339), .B(n2340), .Y(n2337), .VDD(VDD), .GND(VSS) );
NAND2X1 X199 (.A(n2342), .B(n2343), .Y(n2292), .VDD(VDD), .GND(VSS) );
NAND2X1 X200 (.A(n2344), .B(n2345), .Y(n2343), .VDD(VDD), .GND(VSS) );
NAND2X1 X201 (.A(n2349), .B(n2350), .Y(n2341), .VDD(VDD), .GND(VSS) );
NAND2X1 X202 (.A(n2351), .B(n2299), .Y(n2300), .VDD(VDD), .GND(VSS) );
NAND2X1 X203 (.A(n2354), .B(n2355), .Y(n2353), .VDD(VDD), .GND(VSS) );
NAND2X1 X204 (.A(n2356), .B(n2357), .Y(n2354), .VDD(VDD), .GND(VSS) );
NAND2X1 X205 (.A(n2359), .B(n2360), .Y(n2351), .VDD(VDD), .GND(VSS) );
NAND2X1 X206 (.A(N222), .B(N494), .Y(n2312), .VDD(VDD), .GND(VSS) );
NAND2X1 X207 (.A(n2364), .B(n2365), .Y(n2363), .VDD(VDD), .GND(VSS) );
NAND2X1 X208 (.A(n2366), .B(n2364), .Y(n2361), .VDD(VDD), .GND(VSS) );
NAND2X1 X209 (.A(n2367), .B(n2368), .Y(n2364), .VDD(VDD), .GND(VSS) );
NAND2X1 X210 (.A(n2371), .B(N477), .Y(n2370), .VDD(VDD), .GND(VSS) );
NAND2X1 X211 (.A(n2376), .B(n2270), .Y(n2375), .VDD(VDD), .GND(VSS) );
NAND2X1 X212 (.A(N239), .B(n2377), .Y(n2376), .VDD(VDD), .GND(VSS) );
NAND2X1 X213 (.A(n2378), .B(n2379), .Y(n2324), .VDD(VDD), .GND(VSS) );
NAND2X1 X214 (.A(N477), .B(N239), .Y(n2379), .VDD(VDD), .GND(VSS) );
NAND2X1 X215 (.A(N460), .B(N256), .Y(n2326), .VDD(VDD), .GND(VSS) );
NAND2X1 X216 (.A(n2382), .B(n2383), .Y(n2381), .VDD(VDD), .GND(VSS) );
NAND2X1 X217 (.A(N188), .B(N528), .Y(n2294), .VDD(VDD), .GND(VSS) );
NAND2X1 X218 (.A(n2334), .B(n2388), .Y(N6240), .VDD(VDD), .GND(VSS) );
NAND2X1 X219 (.A(n2389), .B(n2390), .Y(n2334), .VDD(VDD), .GND(VSS) );
NAND2X1 X220 (.A(n2391), .B(n2392), .Y(n2390), .VDD(VDD), .GND(VSS) );
NAND2X1 X221 (.A(n2393), .B(n2394), .Y(n2391), .VDD(VDD), .GND(VSS) );
NAND2X1 X222 (.A(n2395), .B(n2396), .Y(n2336), .VDD(VDD), .GND(VSS) );
NAND2X1 X223 (.A(n2397), .B(n2398), .Y(n2395), .VDD(VDD), .GND(VSS) );
NAND2X1 X224 (.A(n2400), .B(n2401), .Y(n2338), .VDD(VDD), .GND(VSS) );
NAND2X1 X225 (.A(n2402), .B(n2403), .Y(n2401), .VDD(VDD), .GND(VSS) );
NAND2X1 X226 (.A(n2407), .B(n2408), .Y(n2399), .VDD(VDD), .GND(VSS) );
NAND2X1 X227 (.A(n2409), .B(n2345), .Y(n2346), .VDD(VDD), .GND(VSS) );
NAND2X1 X228 (.A(n2412), .B(n2413), .Y(n2411), .VDD(VDD), .GND(VSS) );
NAND2X1 X229 (.A(n2417), .B(n2418), .Y(n2409), .VDD(VDD), .GND(VSS) );
NAND2X1 X230 (.A(N205), .B(N494), .Y(n2357), .VDD(VDD), .GND(VSS) );
NAND2X1 X231 (.A(n2422), .B(n2423), .Y(n2421), .VDD(VDD), .GND(VSS) );
NAND2X1 X232 (.A(n2427), .B(n2428), .Y(n2419), .VDD(VDD), .GND(VSS) );
NAND2X1 X233 (.A(N222), .B(N477), .Y(n2368), .VDD(VDD), .GND(VSS) );
NAND2X1 X234 (.A(n2432), .B(n2433), .Y(n2431), .VDD(VDD), .GND(VSS) );
NAND2X1 X235 (.A(n2434), .B(n2432), .Y(n2429), .VDD(VDD), .GND(VSS) );
NAND2X1 X236 (.A(n2435), .B(n2436), .Y(n2432), .VDD(VDD), .GND(VSS) );
NAND2X1 X237 (.A(n2439), .B(N460), .Y(n2438), .VDD(VDD), .GND(VSS) );
NAND2X1 X238 (.A(n2444), .B(n2270), .Y(n2443), .VDD(VDD), .GND(VSS) );
NAND2X1 X239 (.A(N239), .B(n2445), .Y(n2444), .VDD(VDD), .GND(VSS) );
NAND2X1 X240 (.A(n2446), .B(n2447), .Y(n2380), .VDD(VDD), .GND(VSS) );
NAND2X1 X241 (.A(N460), .B(N239), .Y(n2447), .VDD(VDD), .GND(VSS) );
NAND2X1 X242 (.A(N443), .B(N256), .Y(n2382), .VDD(VDD), .GND(VSS) );
NAND2X1 X243 (.A(n2450), .B(n2451), .Y(n2449), .VDD(VDD), .GND(VSS) );
NAND2X1 X244 (.A(N171), .B(N528), .Y(n2340), .VDD(VDD), .GND(VSS) );
NAND2X1 X245 (.A(n2392), .B(n2458), .Y(N6230), .VDD(VDD), .GND(VSS) );
NAND2X1 X246 (.A(n2459), .B(n2460), .Y(n2392), .VDD(VDD), .GND(VSS) );
NAND2X1 X247 (.A(n2461), .B(n2462), .Y(n2460), .VDD(VDD), .GND(VSS) );
NAND2X1 X248 (.A(n2463), .B(n2464), .Y(n2461), .VDD(VDD), .GND(VSS) );
NAND2X1 X249 (.A(n2465), .B(n2466), .Y(n2394), .VDD(VDD), .GND(VSS) );
NAND2X1 X250 (.A(n2467), .B(n2468), .Y(n2465), .VDD(VDD), .GND(VSS) );
NAND2X1 X251 (.A(n2470), .B(n2471), .Y(n2396), .VDD(VDD), .GND(VSS) );
NAND2X1 X252 (.A(n2472), .B(n2473), .Y(n2471), .VDD(VDD), .GND(VSS) );
NAND2X1 X253 (.A(n2477), .B(n2478), .Y(n2469), .VDD(VDD), .GND(VSS) );
NAND2X1 X254 (.A(n2479), .B(n2403), .Y(n2404), .VDD(VDD), .GND(VSS) );
NAND2X1 X255 (.A(n2482), .B(n2483), .Y(n2481), .VDD(VDD), .GND(VSS) );
NAND2X1 X256 (.A(n2487), .B(n2488), .Y(n2479), .VDD(VDD), .GND(VSS) );
NAND2X1 X257 (.A(n2489), .B(n2413), .Y(n2414), .VDD(VDD), .GND(VSS) );
NAND2X1 X258 (.A(n2492), .B(n2493), .Y(n2491), .VDD(VDD), .GND(VSS) );
NAND2X1 X259 (.A(n2497), .B(n2498), .Y(n2489), .VDD(VDD), .GND(VSS) );
NAND2X1 X260 (.A(n2499), .B(n2423), .Y(n2424), .VDD(VDD), .GND(VSS) );
NAND2X1 X261 (.A(n2502), .B(n2503), .Y(n2501), .VDD(VDD), .GND(VSS) );
NAND2X1 X262 (.A(n2504), .B(n2505), .Y(n2502), .VDD(VDD), .GND(VSS) );
NAND2X1 X263 (.A(n2507), .B(n2508), .Y(n2499), .VDD(VDD), .GND(VSS) );
NAND2X1 X264 (.A(N222), .B(N460), .Y(n2436), .VDD(VDD), .GND(VSS) );
NAND2X1 X265 (.A(n2512), .B(n2513), .Y(n2511), .VDD(VDD), .GND(VSS) );
NAND2X1 X266 (.A(n2514), .B(n2512), .Y(n2509), .VDD(VDD), .GND(VSS) );
NAND2X1 X267 (.A(n2515), .B(n2516), .Y(n2512), .VDD(VDD), .GND(VSS) );
NAND2X1 X268 (.A(n2519), .B(N443), .Y(n2518), .VDD(VDD), .GND(VSS) );
NAND2X1 X269 (.A(n2524), .B(n2270), .Y(n2523), .VDD(VDD), .GND(VSS) );
NAND2X1 X270 (.A(N239), .B(n2525), .Y(n2524), .VDD(VDD), .GND(VSS) );
NAND2X1 X271 (.A(n2526), .B(n2527), .Y(n2448), .VDD(VDD), .GND(VSS) );
NAND2X1 X272 (.A(N443), .B(N239), .Y(n2527), .VDD(VDD), .GND(VSS) );
NAND2X1 X273 (.A(N426), .B(N256), .Y(n2450), .VDD(VDD), .GND(VSS) );
NAND2X1 X274 (.A(n2530), .B(n2531), .Y(n2529), .VDD(VDD), .GND(VSS) );
INVX1 X275 (.A(n2202), .AN(n2207), .VDD(VDD), .GND(VSS) );
INVX1 X276 (.A(n2513), .AN(n2517), .VDD(VDD), .GND(VSS) );
XOR2 X277 (.A(n2463), .B(n2464), .Y(n2541), .VDD(VDD), .GND(VSS) );
XOR2 X278 (.A(n2468), .B(n2467), .Y(n2463), .VDD(VDD), .GND(VSS) );
XOR2 X279 (.A(n2475), .B(n2474), .Y(n2552), .VDD(VDD), .GND(VSS) );
XOR2 X280 (.A(n2474), .B(n2558), .Y(n2560), .VDD(VDD), .GND(VSS) );
XOR2 X281 (.A(n2485), .B(n2484), .Y(n2562), .VDD(VDD), .GND(VSS) );
XOR2 X282 (.A(n2484), .B(n2568), .Y(n2570), .VDD(VDD), .GND(VSS) );
XOR2 X283 (.A(n2495), .B(n2494), .Y(n2572), .VDD(VDD), .GND(VSS) );
XOR2 X284 (.A(n2494), .B(n2578), .Y(n2580), .VDD(VDD), .GND(VSS) );
XOR2 X285 (.A(n2505), .B(n2504), .Y(n2582), .VDD(VDD), .GND(VSS) );
XOR2 X286 (.A(n2588), .B(n2505), .Y(n2590), .VDD(VDD), .GND(VSS) );
XOR2 X287 (.A(n2516), .B(n2515), .Y(n2592), .VDD(VDD), .GND(VSS) );
XOR2 X288 (.A(n2598), .B(n2516), .Y(n2600), .VDD(VDD), .GND(VSS) );
XOR2 X289 (.A(n2531), .B(n2530), .Y(n2618), .VDD(VDD), .GND(VSS) );
XOR2 X290 (.A(n2545), .B(n2546), .Y(n2635), .VDD(VDD), .GND(VSS) );
XOR2 X291 (.A(n2550), .B(n2549), .Y(n2545), .VDD(VDD), .GND(VSS) );
XOR2 X292 (.A(n2557), .B(n2556), .Y(n2646), .VDD(VDD), .GND(VSS) );
XOR2 X293 (.A(n2556), .B(n2652), .Y(n2654), .VDD(VDD), .GND(VSS) );
XOR2 X294 (.A(n2567), .B(n2566), .Y(n2656), .VDD(VDD), .GND(VSS) );
XOR2 X295 (.A(n2566), .B(n2662), .Y(n2664), .VDD(VDD), .GND(VSS) );
XOR2 X296 (.A(n2577), .B(n2576), .Y(n2666), .VDD(VDD), .GND(VSS) );
XOR2 X297 (.A(n2576), .B(n2672), .Y(n2674), .VDD(VDD), .GND(VSS) );
XOR2 X298 (.A(n2587), .B(n2586), .Y(n2676), .VDD(VDD), .GND(VSS) );
XOR2 X299 (.A(n2586), .B(n2682), .Y(n2684), .VDD(VDD), .GND(VSS) );
XOR2 X300 (.A(n2597), .B(n2596), .Y(n2686), .VDD(VDD), .GND(VSS) );
XOR2 X301 (.A(n2596), .B(n2692), .Y(n2694), .VDD(VDD), .GND(VSS) );
XOR2 X302 (.A(n2608), .B(n2607), .Y(n2696), .VDD(VDD), .GND(VSS) );
XOR2 X303 (.A(n2702), .B(n2608), .Y(n2704), .VDD(VDD), .GND(VSS) );
XOR2 X304 (.A(n2623), .B(n2622), .Y(n2722), .VDD(VDD), .GND(VSS) );
XOR2 X305 (.A(n2639), .B(n2640), .Y(n2741), .VDD(VDD), .GND(VSS) );
XOR2 X306 (.A(n2644), .B(n2643), .Y(n2639), .VDD(VDD), .GND(VSS) );
XOR2 X307 (.A(n2651), .B(n2650), .Y(n2752), .VDD(VDD), .GND(VSS) );
XOR2 X308 (.A(n2650), .B(n2758), .Y(n2760), .VDD(VDD), .GND(VSS) );
XOR2 X309 (.A(n2661), .B(n2660), .Y(n2762), .VDD(VDD), .GND(VSS) );
XOR2 X310 (.A(n2660), .B(n2768), .Y(n2770), .VDD(VDD), .GND(VSS) );
XOR2 X311 (.A(n2671), .B(n2670), .Y(n2772), .VDD(VDD), .GND(VSS) );
XOR2 X312 (.A(n2670), .B(n2778), .Y(n2780), .VDD(VDD), .GND(VSS) );
XOR2 X313 (.A(n2681), .B(n2680), .Y(n2782), .VDD(VDD), .GND(VSS) );
XOR2 X314 (.A(n2680), .B(n2788), .Y(n2790), .VDD(VDD), .GND(VSS) );
XOR2 X315 (.A(n2691), .B(n2690), .Y(n2792), .VDD(VDD), .GND(VSS) );
XOR2 X316 (.A(n2690), .B(n2798), .Y(n2800), .VDD(VDD), .GND(VSS) );
XOR2 X317 (.A(n2701), .B(n2700), .Y(n2802), .VDD(VDD), .GND(VSS) );
XOR2 X318 (.A(n2808), .B(n2701), .Y(n2810), .VDD(VDD), .GND(VSS) );
XOR2 X319 (.A(n2712), .B(n2711), .Y(n2812), .VDD(VDD), .GND(VSS) );
XOR2 X320 (.A(n2818), .B(n2712), .Y(n2820), .VDD(VDD), .GND(VSS) );
OR2X1 X321 (.A(n2541), .B(n2542), .VDD(VDD), .VSS(VSS), .Y(n2540) );
OR2X1 X322 (.A(n2556), .B(n2557), .VDD(VDD), .VSS(VSS), .Y(n2554) );
OR2X1 X323 (.A(n2566), .B(n2567), .VDD(VDD), .VSS(VSS), .Y(n2564) );
OR2X1 X324 (.A(n2576), .B(n2577), .VDD(VDD), .VSS(VSS), .Y(n2574) );
OR2X1 X325 (.A(n2586), .B(n2587), .VDD(VDD), .VSS(VSS), .Y(n2584) );
OR2X1 X326 (.A(n2596), .B(n2597), .VDD(VDD), .VSS(VSS), .Y(n2594) );
OR2X1 X327 (.A(n2635), .B(n2636), .VDD(VDD), .VSS(VSS), .Y(n2634) );
OR2X1 X328 (.A(n2650), .B(n2651), .VDD(VDD), .VSS(VSS), .Y(n2648) );
OR2X1 X329 (.A(n2660), .B(n2661), .VDD(VDD), .VSS(VSS), .Y(n2658) );
OR2X1 X330 (.A(n2670), .B(n2671), .VDD(VDD), .VSS(VSS), .Y(n2668) );
OR2X1 X331 (.A(n2680), .B(n2681), .VDD(VDD), .VSS(VSS), .Y(n2678) );
OR2X1 X332 (.A(n2690), .B(n2691), .VDD(VDD), .VSS(VSS), .Y(n2688) );
OR2X1 X333 (.A(n2741), .B(n2742), .VDD(VDD), .VSS(VSS), .Y(n2740) );
OR2X1 X334 (.A(n2756), .B(n2757), .VDD(VDD), .VSS(VSS), .Y(n2754) );
OR2X1 X335 (.A(n2766), .B(n2767), .VDD(VDD), .VSS(VSS), .Y(n2764) );
OR2X1 X336 (.A(n2776), .B(n2777), .VDD(VDD), .VSS(VSS), .Y(n2774) );
OR2X1 X337 (.A(n2786), .B(n2787), .VDD(VDD), .VSS(VSS), .Y(n2784) );
OR2X1 X338 (.A(n2796), .B(n2797), .VDD(VDD), .VSS(VSS), .Y(n2794) );
OR2X1 X339 (.A(n2806), .B(n2807), .VDD(VDD), .VSS(VSS), .Y(n2804) );
OR2X1 X340 (.A(n2816), .B(n2817), .VDD(VDD), .VSS(VSS), .Y(n2814) );
AND2X1 X341 (.A(n2593), .B(n2592), .VDD(VDD), .VSS(VSS), .Y(n2532) );
AND2X1 X342 (.A(n2583), .B(n2582), .VDD(VDD), .VSS(VSS), .Y(n2534) );
AND2X1 X343 (.A(n2573), .B(n2572), .VDD(VDD), .VSS(VSS), .Y(n2536) );
AND2X1 X344 (.A(n2563), .B(n2562), .VDD(VDD), .VSS(VSS), .Y(n2538) );
AND2X1 X345 (.A(n2551), .B(n2466), .VDD(VDD), .VSS(VSS), .Y(n2467) );
AND2X1 X346 (.A(N511), .B(N154), .VDD(VDD), .VSS(VSS), .Y(n2475) );
AND2X1 X347 (.A(N494), .B(N171), .VDD(VDD), .VSS(VSS), .Y(n2485) );
AND2X1 X348 (.A(N477), .B(N188), .VDD(VDD), .VSS(VSS), .Y(n2495) );
AND2X1 X349 (.A(n2503), .B(n2591), .VDD(VDD), .VSS(VSS), .Y(n2504) );
AND2X1 X350 (.A(n2513), .B(n2601), .VDD(VDD), .VSS(VSS), .Y(n2515) );
AND2X1 X351 (.A(n2528), .B(n2610), .VDD(VDD), .VSS(VSS), .Y(n2602) );
AND2X1 X352 (.A(n2621), .B(n2620), .VDD(VDD), .VSS(VSS), .Y(n2614) );
AND2X1 X353 (.A(n2707), .B(n2706), .VDD(VDD), .VSS(VSS), .Y(n2609) );
AND2X1 X354 (.A(n2697), .B(n2696), .VDD(VDD), .VSS(VSS), .Y(n2624) );
AND2X1 X355 (.A(n2687), .B(n2686), .VDD(VDD), .VSS(VSS), .Y(n2626) );
AND2X1 X356 (.A(n2677), .B(n2676), .VDD(VDD), .VSS(VSS), .Y(n2628) );
AND2X1 X357 (.A(n2667), .B(n2666), .VDD(VDD), .VSS(VSS), .Y(n2630) );
AND2X1 X358 (.A(n2657), .B(n2656), .VDD(VDD), .VSS(VSS), .Y(n2632) );
AND2X1 X359 (.A(n2645), .B(n2548), .VDD(VDD), .VSS(VSS), .Y(n2549) );
AND2X1 X360 (.A(N511), .B(N137), .VDD(VDD), .VSS(VSS), .Y(n2557) );
AND2X1 X361 (.A(N494), .B(N154), .VDD(VDD), .VSS(VSS), .Y(n2567) );
AND2X1 X362 (.A(N477), .B(N171), .VDD(VDD), .VSS(VSS), .Y(n2577) );
AND2X1 X363 (.A(N460), .B(N188), .VDD(VDD), .VSS(VSS), .Y(n2587) );
AND2X1 X364 (.A(N443), .B(N205), .VDD(VDD), .VSS(VSS), .Y(n2597) );
AND2X1 X365 (.A(n2605), .B(n2705), .VDD(VDD), .VSS(VSS), .Y(n2607) );
AND2X1 X366 (.A(n2620), .B(n2714), .VDD(VDD), .VSS(VSS), .Y(n2706) );
AND2X1 X367 (.A(n2725), .B(n2724), .VDD(VDD), .VSS(VSS), .Y(n2718) );
AND2X1 X368 (.A(n2823), .B(n2822), .VDD(VDD), .VSS(VSS), .Y(n2713) );
AND2X1 X369 (.A(n2701), .B(n2700), .VDD(VDD), .VSS(VSS), .Y(n2729) );
AND2X1 X370 (.A(n2813), .B(n2812), .VDD(VDD), .VSS(VSS), .Y(n2728) );
AND2X1 X371 (.A(n2803), .B(n2802), .VDD(VDD), .VSS(VSS), .Y(n2730) );
AND2X1 X372 (.A(n2793), .B(n2792), .VDD(VDD), .VSS(VSS), .Y(n2732) );
AND2X1 X373 (.A(n2783), .B(n2782), .VDD(VDD), .VSS(VSS), .Y(n2734) );
AND2X1 X374 (.A(n2773), .B(n2772), .VDD(VDD), .VSS(VSS), .Y(n2736) );
AND2X1 X375 (.A(n2763), .B(n2762), .VDD(VDD), .VSS(VSS), .Y(n2738) );
AND2X1 X376 (.A(n2751), .B(n2642), .VDD(VDD), .VSS(VSS), .Y(n2643) );
AND2X1 X377 (.A(N511), .B(N120), .VDD(VDD), .VSS(VSS), .Y(n2651) );
AND2X1 X378 (.A(N494), .B(N137), .VDD(VDD), .VSS(VSS), .Y(n2661) );
AND2X1 X379 (.A(N477), .B(N154), .VDD(VDD), .VSS(VSS), .Y(n2671) );
AND2X1 X380 (.A(N460), .B(N171), .VDD(VDD), .VSS(VSS), .Y(n2681) );
AND2X1 X381 (.A(N443), .B(N188), .VDD(VDD), .VSS(VSS), .Y(n2691) );
AND2X1 X382 (.A(n2699), .B(n2811), .VDD(VDD), .VSS(VSS), .Y(n2700) );
AND2X1 X383 (.A(n2709), .B(n2821), .VDD(VDD), .VSS(VSS), .Y(n2711) );
AND2X1 X384 (.A(n2724), .B(n2830), .VDD(VDD), .VSS(VSS), .Y(n2822) );
NOR2X1 X385 (.A(n2534), .B(n2535), .Y(n2497), .VDD(VDD), .GND(VSS) );
NOR2X1 X386 (.A(n2495), .B(n2494), .Y(n2535), .VDD(VDD), .GND(VSS) );
NOR2X1 X387 (.A(n2536), .B(n2537), .Y(n2487), .VDD(VDD), .GND(VSS) );
NOR2X1 X388 (.A(n2485), .B(n2484), .Y(n2537), .VDD(VDD), .GND(VSS) );
NOR2X1 X389 (.A(n2538), .B(n2539), .Y(n2477), .VDD(VDD), .GND(VSS) );
NOR2X1 X390 (.A(n2475), .B(n2474), .Y(n2539), .VDD(VDD), .GND(VSS) );
NOR2X1 X391 (.A(n2609), .B(n2602), .Y(n2606), .VDD(VDD), .GND(VSS) );
NOR2X1 X392 (.A(n2612), .B(n2613), .Y(n2611), .VDD(VDD), .GND(VSS) );
NOR2X1 X393 (.A(n2614), .B(n2615), .Y(n2613), .VDD(VDD), .GND(VSS) );
NOR2X1 X394 (.A(N409), .B(n2531), .Y(n2612), .VDD(VDD), .GND(VSS) );
NOR2X1 X395 (.A(n2624), .B(n2625), .Y(n2599), .VDD(VDD), .GND(VSS) );
NOR2X1 X396 (.A(n2597), .B(n2596), .Y(n2625), .VDD(VDD), .GND(VSS) );
NOR2X1 X397 (.A(n2626), .B(n2627), .Y(n2589), .VDD(VDD), .GND(VSS) );
NOR2X1 X398 (.A(n2587), .B(n2586), .Y(n2627), .VDD(VDD), .GND(VSS) );
NOR2X1 X399 (.A(n2628), .B(n2629), .Y(n2579), .VDD(VDD), .GND(VSS) );
NOR2X1 X400 (.A(n2577), .B(n2576), .Y(n2629), .VDD(VDD), .GND(VSS) );
NOR2X1 X401 (.A(n2630), .B(n2631), .Y(n2569), .VDD(VDD), .GND(VSS) );
NOR2X1 X402 (.A(n2567), .B(n2566), .Y(n2631), .VDD(VDD), .GND(VSS) );
NOR2X1 X403 (.A(n2632), .B(n2633), .Y(n2559), .VDD(VDD), .GND(VSS) );
NOR2X1 X404 (.A(n2557), .B(n2556), .Y(n2633), .VDD(VDD), .GND(VSS) );
NOR2X1 X405 (.A(n2713), .B(n2706), .Y(n2710), .VDD(VDD), .GND(VSS) );
NOR2X1 X406 (.A(n2716), .B(n2717), .Y(n2715), .VDD(VDD), .GND(VSS) );
NOR2X1 X407 (.A(n2718), .B(n2719), .Y(n2717), .VDD(VDD), .GND(VSS) );
NOR2X1 X408 (.A(N392), .B(n2623), .Y(n2716), .VDD(VDD), .GND(VSS) );
NOR2X1 X409 (.A(n2728), .B(n2729), .Y(n2703), .VDD(VDD), .GND(VSS) );
NOR2X1 X410 (.A(n2730), .B(n2731), .Y(n2693), .VDD(VDD), .GND(VSS) );
NOR2X1 X411 (.A(n2691), .B(n2690), .Y(n2731), .VDD(VDD), .GND(VSS) );
NOR2X1 X412 (.A(n2732), .B(n2733), .Y(n2683), .VDD(VDD), .GND(VSS) );
NOR2X1 X413 (.A(n2681), .B(n2680), .Y(n2733), .VDD(VDD), .GND(VSS) );
NOR2X1 X414 (.A(n2734), .B(n2735), .Y(n2673), .VDD(VDD), .GND(VSS) );
NOR2X1 X415 (.A(n2671), .B(n2670), .Y(n2735), .VDD(VDD), .GND(VSS) );
NOR2X1 X416 (.A(n2736), .B(n2737), .Y(n2663), .VDD(VDD), .GND(VSS) );
NOR2X1 X417 (.A(n2661), .B(n2660), .Y(n2737), .VDD(VDD), .GND(VSS) );
NOR2X1 X418 (.A(n2738), .B(n2739), .Y(n2653), .VDD(VDD), .GND(VSS) );
NOR2X1 X419 (.A(n2651), .B(n2650), .Y(n2739), .VDD(VDD), .GND(VSS) );
NOR2X1 X420 (.A(n2829), .B(n2822), .Y(n2826), .VDD(VDD), .GND(VSS) );
NOR2X1 X421 (.A(n2832), .B(n2833), .Y(n2831), .VDD(VDD), .GND(VSS) );
NOR2X1 X422 (.A(n2834), .B(n2835), .Y(n2833), .VDD(VDD), .GND(VSS) );
NOR2X1 X423 (.A(N375), .B(n2727), .Y(n2832), .VDD(VDD), .GND(VSS) );
NAND2X1 X424 (.A(N154), .B(N528), .Y(n2398), .VDD(VDD), .GND(VSS) );
NAND2X1 X425 (.A(n2462), .B(n2540), .Y(N6220), .VDD(VDD), .GND(VSS) );
NAND2X1 X426 (.A(n2541), .B(n2542), .Y(n2462), .VDD(VDD), .GND(VSS) );
NAND2X1 X427 (.A(n2543), .B(n2544), .Y(n2542), .VDD(VDD), .GND(VSS) );
NAND2X1 X428 (.A(n2545), .B(n2546), .Y(n2543), .VDD(VDD), .GND(VSS) );
NAND2X1 X429 (.A(n2547), .B(n2548), .Y(n2464), .VDD(VDD), .GND(VSS) );
NAND2X1 X430 (.A(n2549), .B(n2550), .Y(n2547), .VDD(VDD), .GND(VSS) );
NAND2X1 X431 (.A(n2552), .B(n2553), .Y(n2466), .VDD(VDD), .GND(VSS) );
NAND2X1 X432 (.A(n2554), .B(n2555), .Y(n2553), .VDD(VDD), .GND(VSS) );
NAND2X1 X433 (.A(n2559), .B(n2560), .Y(n2551), .VDD(VDD), .GND(VSS) );
NAND2X1 X434 (.A(n2561), .B(n2473), .Y(n2474), .VDD(VDD), .GND(VSS) );
NAND2X1 X435 (.A(n2564), .B(n2565), .Y(n2563), .VDD(VDD), .GND(VSS) );
NAND2X1 X436 (.A(n2569), .B(n2570), .Y(n2561), .VDD(VDD), .GND(VSS) );
NAND2X1 X437 (.A(n2571), .B(n2483), .Y(n2484), .VDD(VDD), .GND(VSS) );
NAND2X1 X438 (.A(n2574), .B(n2575), .Y(n2573), .VDD(VDD), .GND(VSS) );
NAND2X1 X439 (.A(n2579), .B(n2580), .Y(n2571), .VDD(VDD), .GND(VSS) );
NAND2X1 X440 (.A(n2581), .B(n2493), .Y(n2494), .VDD(VDD), .GND(VSS) );
NAND2X1 X441 (.A(n2584), .B(n2585), .Y(n2583), .VDD(VDD), .GND(VSS) );
NAND2X1 X442 (.A(n2589), .B(n2590), .Y(n2581), .VDD(VDD), .GND(VSS) );
NAND2X1 X443 (.A(N205), .B(N460), .Y(n2505), .VDD(VDD), .GND(VSS) );
NAND2X1 X444 (.A(n2594), .B(n2595), .Y(n2593), .VDD(VDD), .GND(VSS) );
NAND2X1 X445 (.A(n2599), .B(n2600), .Y(n2591), .VDD(VDD), .GND(VSS) );
NAND2X1 X446 (.A(N222), .B(N443), .Y(n2516), .VDD(VDD), .GND(VSS) );
NAND2X1 X447 (.A(n2602), .B(n2603), .Y(n2513), .VDD(VDD), .GND(VSS) );
NAND2X1 X448 (.A(n2604), .B(n2605), .Y(n2603), .VDD(VDD), .GND(VSS) );
NAND2X1 X449 (.A(n2606), .B(n2604), .Y(n2601), .VDD(VDD), .GND(VSS) );
NAND2X1 X450 (.A(n2607), .B(n2608), .Y(n2604), .VDD(VDD), .GND(VSS) );
NAND2X1 X451 (.A(n2611), .B(N426), .Y(n2610), .VDD(VDD), .GND(VSS) );
NAND2X1 X452 (.A(n2616), .B(n2270), .Y(n2615), .VDD(VDD), .GND(VSS) );
NAND2X1 X453 (.A(N239), .B(n2617), .Y(n2616), .VDD(VDD), .GND(VSS) );
NAND2X1 X454 (.A(n2618), .B(n2619), .Y(n2528), .VDD(VDD), .GND(VSS) );
NAND2X1 X455 (.A(N426), .B(N239), .Y(n2619), .VDD(VDD), .GND(VSS) );
NAND2X1 X456 (.A(N409), .B(N256), .Y(n2530), .VDD(VDD), .GND(VSS) );
NAND2X1 X457 (.A(n2622), .B(n2623), .Y(n2621), .VDD(VDD), .GND(VSS) );
NAND2X1 X458 (.A(N137), .B(N528), .Y(n2468), .VDD(VDD), .GND(VSS) );
NAND2X1 X459 (.A(n2544), .B(n2634), .Y(N6210), .VDD(VDD), .GND(VSS) );
NAND2X1 X460 (.A(n2635), .B(n2636), .Y(n2544), .VDD(VDD), .GND(VSS) );
NAND2X1 X461 (.A(n2637), .B(n2638), .Y(n2636), .VDD(VDD), .GND(VSS) );
NAND2X1 X462 (.A(n2639), .B(n2640), .Y(n2637), .VDD(VDD), .GND(VSS) );
NAND2X1 X463 (.A(n2641), .B(n2642), .Y(n2546), .VDD(VDD), .GND(VSS) );
NAND2X1 X464 (.A(n2643), .B(n2644), .Y(n2641), .VDD(VDD), .GND(VSS) );
NAND2X1 X465 (.A(n2646), .B(n2647), .Y(n2548), .VDD(VDD), .GND(VSS) );
NAND2X1 X466 (.A(n2648), .B(n2649), .Y(n2647), .VDD(VDD), .GND(VSS) );
NAND2X1 X467 (.A(n2653), .B(n2654), .Y(n2645), .VDD(VDD), .GND(VSS) );
NAND2X1 X468 (.A(n2655), .B(n2555), .Y(n2556), .VDD(VDD), .GND(VSS) );
NAND2X1 X469 (.A(n2658), .B(n2659), .Y(n2657), .VDD(VDD), .GND(VSS) );
NAND2X1 X470 (.A(n2663), .B(n2664), .Y(n2655), .VDD(VDD), .GND(VSS) );
NAND2X1 X471 (.A(n2665), .B(n2565), .Y(n2566), .VDD(VDD), .GND(VSS) );
NAND2X1 X472 (.A(n2668), .B(n2669), .Y(n2667), .VDD(VDD), .GND(VSS) );
NAND2X1 X473 (.A(n2673), .B(n2674), .Y(n2665), .VDD(VDD), .GND(VSS) );
NAND2X1 X474 (.A(n2675), .B(n2575), .Y(n2576), .VDD(VDD), .GND(VSS) );
NAND2X1 X475 (.A(n2678), .B(n2679), .Y(n2677), .VDD(VDD), .GND(VSS) );
NAND2X1 X476 (.A(n2683), .B(n2684), .Y(n2675), .VDD(VDD), .GND(VSS) );
NAND2X1 X477 (.A(n2685), .B(n2585), .Y(n2586), .VDD(VDD), .GND(VSS) );
NAND2X1 X478 (.A(n2688), .B(n2689), .Y(n2687), .VDD(VDD), .GND(VSS) );
NAND2X1 X479 (.A(n2693), .B(n2694), .Y(n2685), .VDD(VDD), .GND(VSS) );
NAND2X1 X480 (.A(n2695), .B(n2595), .Y(n2596), .VDD(VDD), .GND(VSS) );
NAND2X1 X481 (.A(n2698), .B(n2699), .Y(n2697), .VDD(VDD), .GND(VSS) );
NAND2X1 X482 (.A(n2700), .B(n2701), .Y(n2698), .VDD(VDD), .GND(VSS) );
NAND2X1 X483 (.A(n2703), .B(n2704), .Y(n2695), .VDD(VDD), .GND(VSS) );
NAND2X1 X484 (.A(N222), .B(N426), .Y(n2608), .VDD(VDD), .GND(VSS) );
NAND2X1 X485 (.A(n2708), .B(n2709), .Y(n2707), .VDD(VDD), .GND(VSS) );
NAND2X1 X486 (.A(n2710), .B(n2708), .Y(n2705), .VDD(VDD), .GND(VSS) );
NAND2X1 X487 (.A(n2711), .B(n2712), .Y(n2708), .VDD(VDD), .GND(VSS) );
NAND2X1 X488 (.A(n2715), .B(N409), .Y(n2714), .VDD(VDD), .GND(VSS) );
NAND2X1 X489 (.A(n2720), .B(n2270), .Y(n2719), .VDD(VDD), .GND(VSS) );
NAND2X1 X490 (.A(N239), .B(n2721), .Y(n2720), .VDD(VDD), .GND(VSS) );
NAND2X1 X491 (.A(n2722), .B(n2723), .Y(n2620), .VDD(VDD), .GND(VSS) );
NAND2X1 X492 (.A(N409), .B(N239), .Y(n2723), .VDD(VDD), .GND(VSS) );
NAND2X1 X493 (.A(N392), .B(N256), .Y(n2622), .VDD(VDD), .GND(VSS) );
NAND2X1 X494 (.A(n2726), .B(n2727), .Y(n2725), .VDD(VDD), .GND(VSS) );
NAND2X1 X495 (.A(N120), .B(N528), .Y(n2550), .VDD(VDD), .GND(VSS) );
NAND2X1 X496 (.A(n2638), .B(n2740), .Y(N6200), .VDD(VDD), .GND(VSS) );
NAND2X1 X497 (.A(n2741), .B(n2742), .Y(n2638), .VDD(VDD), .GND(VSS) );
NAND2X1 X498 (.A(n2743), .B(n2744), .Y(n2742), .VDD(VDD), .GND(VSS) );
NAND2X1 X499 (.A(n2745), .B(n2746), .Y(n2743), .VDD(VDD), .GND(VSS) );
NAND2X1 X500 (.A(n2747), .B(n2748), .Y(n2640), .VDD(VDD), .GND(VSS) );
NAND2X1 X501 (.A(n2749), .B(n2750), .Y(n2747), .VDD(VDD), .GND(VSS) );
NAND2X1 X502 (.A(n2752), .B(n2753), .Y(n2642), .VDD(VDD), .GND(VSS) );
NAND2X1 X503 (.A(n2754), .B(n2755), .Y(n2753), .VDD(VDD), .GND(VSS) );
NAND2X1 X504 (.A(n2759), .B(n2760), .Y(n2751), .VDD(VDD), .GND(VSS) );
NAND2X1 X505 (.A(n2761), .B(n2649), .Y(n2650), .VDD(VDD), .GND(VSS) );
NAND2X1 X506 (.A(n2764), .B(n2765), .Y(n2763), .VDD(VDD), .GND(VSS) );
NAND2X1 X507 (.A(n2769), .B(n2770), .Y(n2761), .VDD(VDD), .GND(VSS) );
NAND2X1 X508 (.A(n2771), .B(n2659), .Y(n2660), .VDD(VDD), .GND(VSS) );
NAND2X1 X509 (.A(n2774), .B(n2775), .Y(n2773), .VDD(VDD), .GND(VSS) );
NAND2X1 X510 (.A(n2779), .B(n2780), .Y(n2771), .VDD(VDD), .GND(VSS) );
NAND2X1 X511 (.A(n2781), .B(n2669), .Y(n2670), .VDD(VDD), .GND(VSS) );
NAND2X1 X512 (.A(n2784), .B(n2785), .Y(n2783), .VDD(VDD), .GND(VSS) );
NAND2X1 X513 (.A(n2789), .B(n2790), .Y(n2781), .VDD(VDD), .GND(VSS) );
NAND2X1 X514 (.A(n2791), .B(n2679), .Y(n2680), .VDD(VDD), .GND(VSS) );
NAND2X1 X515 (.A(n2794), .B(n2795), .Y(n2793), .VDD(VDD), .GND(VSS) );
NAND2X1 X516 (.A(n2799), .B(n2800), .Y(n2791), .VDD(VDD), .GND(VSS) );
NAND2X1 X517 (.A(n2801), .B(n2689), .Y(n2690), .VDD(VDD), .GND(VSS) );
NAND2X1 X518 (.A(n2804), .B(n2805), .Y(n2803), .VDD(VDD), .GND(VSS) );
NAND2X1 X519 (.A(n2809), .B(n2810), .Y(n2801), .VDD(VDD), .GND(VSS) );
NAND2X1 X520 (.A(N205), .B(N426), .Y(n2701), .VDD(VDD), .GND(VSS) );
NAND2X1 X521 (.A(n2814), .B(n2815), .Y(n2813), .VDD(VDD), .GND(VSS) );
NAND2X1 X522 (.A(n2819), .B(n2820), .Y(n2811), .VDD(VDD), .GND(VSS) );
NAND2X1 X523 (.A(N222), .B(N409), .Y(n2712), .VDD(VDD), .GND(VSS) );
NAND2X1 X524 (.A(n2824), .B(n2825), .Y(n2823), .VDD(VDD), .GND(VSS) );
NAND2X1 X525 (.A(n2826), .B(n2824), .Y(n2821), .VDD(VDD), .GND(VSS) );
NAND2X1 X526 (.A(n2827), .B(n2828), .Y(n2824), .VDD(VDD), .GND(VSS) );
NAND2X1 X527 (.A(n2831), .B(N392), .Y(n2830), .VDD(VDD), .GND(VSS) );
NAND2X1 X528 (.A(n2836), .B(n2270), .Y(n2835), .VDD(VDD), .GND(VSS) );
NAND2X1 X529 (.A(N239), .B(n2837), .Y(n2836), .VDD(VDD), .GND(VSS) );
INVX1 X530 (.A(n2727), .AN(n2834), .VDD(VDD), .GND(VSS) );
XOR2 X531 (.A(n2727), .B(n2726), .Y(n2838), .VDD(VDD), .GND(VSS) );
XOR2 X532 (.A(n2745), .B(n2746), .Y(n2859), .VDD(VDD), .GND(VSS) );
XOR2 X533 (.A(n2750), .B(n2749), .Y(n2745), .VDD(VDD), .GND(VSS) );
XOR2 X534 (.A(n2757), .B(n2756), .Y(n2870), .VDD(VDD), .GND(VSS) );
XOR2 X535 (.A(n2756), .B(n2876), .Y(n2878), .VDD(VDD), .GND(VSS) );
XOR2 X536 (.A(n2767), .B(n2766), .Y(n2880), .VDD(VDD), .GND(VSS) );
XOR2 X537 (.A(n2766), .B(n2886), .Y(n2888), .VDD(VDD), .GND(VSS) );
XOR2 X538 (.A(n2777), .B(n2776), .Y(n2890), .VDD(VDD), .GND(VSS) );
XOR2 X539 (.A(n2776), .B(n2896), .Y(n2898), .VDD(VDD), .GND(VSS) );
XOR2 X540 (.A(n2787), .B(n2786), .Y(n2900), .VDD(VDD), .GND(VSS) );
XOR2 X541 (.A(n2786), .B(n2906), .Y(n2908), .VDD(VDD), .GND(VSS) );
XOR2 X542 (.A(n2797), .B(n2796), .Y(n2910), .VDD(VDD), .GND(VSS) );
XOR2 X543 (.A(n2796), .B(n2916), .Y(n2918), .VDD(VDD), .GND(VSS) );
XOR2 X544 (.A(n2807), .B(n2806), .Y(n2920), .VDD(VDD), .GND(VSS) );
XOR2 X545 (.A(n2806), .B(n2926), .Y(n2928), .VDD(VDD), .GND(VSS) );
XOR2 X546 (.A(n2817), .B(n2816), .Y(n2930), .VDD(VDD), .GND(VSS) );
XOR2 X547 (.A(n2816), .B(n2936), .Y(n2938), .VDD(VDD), .GND(VSS) );
XOR2 X548 (.A(n2828), .B(n2827), .Y(n2940), .VDD(VDD), .GND(VSS) );
XOR2 X549 (.A(n2946), .B(n2828), .Y(n2948), .VDD(VDD), .GND(VSS) );
XOR2 X550 (.A(n2843), .B(n2842), .Y(n2966), .VDD(VDD), .GND(VSS) );
XOR2 X551 (.A(n2863), .B(n2864), .Y(n2989), .VDD(VDD), .GND(VSS) );
XOR2 X552 (.A(n2868), .B(n2867), .Y(n2863), .VDD(VDD), .GND(VSS) );
XOR2 X553 (.A(n2875), .B(n2874), .Y(n3000), .VDD(VDD), .GND(VSS) );
XOR2 X554 (.A(n2874), .B(n3006), .Y(n3008), .VDD(VDD), .GND(VSS) );
XOR2 X555 (.A(n2885), .B(n2884), .Y(n3010), .VDD(VDD), .GND(VSS) );
XOR2 X556 (.A(n2884), .B(n3016), .Y(n3018), .VDD(VDD), .GND(VSS) );
XOR2 X557 (.A(n2895), .B(n2894), .Y(n3020), .VDD(VDD), .GND(VSS) );
XOR2 X558 (.A(n2894), .B(n3026), .Y(n3028), .VDD(VDD), .GND(VSS) );
XOR2 X559 (.A(n2905), .B(n2904), .Y(n3030), .VDD(VDD), .GND(VSS) );
XOR2 X560 (.A(n2904), .B(n3036), .Y(n3038), .VDD(VDD), .GND(VSS) );
XOR2 X561 (.A(n2915), .B(n2914), .Y(n3040), .VDD(VDD), .GND(VSS) );
XOR2 X562 (.A(n2914), .B(n3046), .Y(n3048), .VDD(VDD), .GND(VSS) );
XOR2 X563 (.A(n2925), .B(n2924), .Y(n3050), .VDD(VDD), .GND(VSS) );
XOR2 X564 (.A(n2924), .B(n3056), .Y(n3058), .VDD(VDD), .GND(VSS) );
XOR2 X565 (.A(n2935), .B(n2934), .Y(n3060), .VDD(VDD), .GND(VSS) );
XOR2 X566 (.A(n2934), .B(n3066), .Y(n3068), .VDD(VDD), .GND(VSS) );
XOR2 X567 (.A(n2945), .B(n2944), .Y(n3070), .VDD(VDD), .GND(VSS) );
XOR2 X568 (.A(n3076), .B(n2945), .Y(n3078), .VDD(VDD), .GND(VSS) );
XOR2 X569 (.A(n2956), .B(n2955), .Y(n3080), .VDD(VDD), .GND(VSS) );
XOR2 X570 (.A(n3086), .B(n2956), .Y(n3088), .VDD(VDD), .GND(VSS) );
XOR2 X571 (.A(n2971), .B(n2970), .Y(n3106), .VDD(VDD), .GND(VSS) );
XOR2 X572 (.A(n2993), .B(n2994), .Y(n3131), .VDD(VDD), .GND(VSS) );
OR2X1 X573 (.A(n2859), .B(n2860), .VDD(VDD), .VSS(VSS), .Y(n2858) );
OR2X1 X574 (.A(n2874), .B(n2875), .VDD(VDD), .VSS(VSS), .Y(n2872) );
OR2X1 X575 (.A(n2884), .B(n2885), .VDD(VDD), .VSS(VSS), .Y(n2882) );
OR2X1 X576 (.A(n2894), .B(n2895), .VDD(VDD), .VSS(VSS), .Y(n2892) );
OR2X1 X577 (.A(n2904), .B(n2905), .VDD(VDD), .VSS(VSS), .Y(n2902) );
OR2X1 X578 (.A(n2914), .B(n2915), .VDD(VDD), .VSS(VSS), .Y(n2912) );
OR2X1 X579 (.A(n2924), .B(n2925), .VDD(VDD), .VSS(VSS), .Y(n2922) );
OR2X1 X580 (.A(n2934), .B(n2935), .VDD(VDD), .VSS(VSS), .Y(n2932) );
OR2X1 X581 (.A(n2989), .B(n2990), .VDD(VDD), .VSS(VSS), .Y(n2988) );
OR2X1 X582 (.A(n3004), .B(n3005), .VDD(VDD), .VSS(VSS), .Y(n3002) );
OR2X1 X583 (.A(n3014), .B(n3015), .VDD(VDD), .VSS(VSS), .Y(n3012) );
OR2X1 X584 (.A(n3024), .B(n3025), .VDD(VDD), .VSS(VSS), .Y(n3022) );
OR2X1 X585 (.A(n3034), .B(n3035), .VDD(VDD), .VSS(VSS), .Y(n3032) );
OR2X1 X586 (.A(n3044), .B(n3045), .VDD(VDD), .VSS(VSS), .Y(n3042) );
OR2X1 X587 (.A(n3054), .B(n3055), .VDD(VDD), .VSS(VSS), .Y(n3052) );
OR2X1 X588 (.A(n3064), .B(n3065), .VDD(VDD), .VSS(VSS), .Y(n3062) );
OR2X1 X589 (.A(n3074), .B(n3075), .VDD(VDD), .VSS(VSS), .Y(n3072) );
OR2X1 X590 (.A(n3084), .B(n3085), .VDD(VDD), .VSS(VSS), .Y(n3082) );
OR2X1 X591 (.A(n3131), .B(n3132), .VDD(VDD), .VSS(VSS), .Y(n3130) );
AND2X1 X592 (.A(n2951), .B(n2950), .VDD(VDD), .VSS(VSS), .Y(n2829) );
AND2X1 X593 (.A(n2941), .B(n2940), .VDD(VDD), .VSS(VSS), .Y(n2844) );
AND2X1 X594 (.A(n2931), .B(n2930), .VDD(VDD), .VSS(VSS), .Y(n2846) );
AND2X1 X595 (.A(n2921), .B(n2920), .VDD(VDD), .VSS(VSS), .Y(n2848) );
AND2X1 X596 (.A(n2911), .B(n2910), .VDD(VDD), .VSS(VSS), .Y(n2850) );
AND2X1 X597 (.A(n2901), .B(n2900), .VDD(VDD), .VSS(VSS), .Y(n2852) );
AND2X1 X598 (.A(n2891), .B(n2890), .VDD(VDD), .VSS(VSS), .Y(n2854) );
AND2X1 X599 (.A(n2881), .B(n2880), .VDD(VDD), .VSS(VSS), .Y(n2856) );
AND2X1 X600 (.A(n2869), .B(n2748), .VDD(VDD), .VSS(VSS), .Y(n2749) );
AND2X1 X601 (.A(N511), .B(N103), .VDD(VDD), .VSS(VSS), .Y(n2757) );
AND2X1 X602 (.A(N494), .B(N120), .VDD(VDD), .VSS(VSS), .Y(n2767) );
AND2X1 X603 (.A(N477), .B(N137), .VDD(VDD), .VSS(VSS), .Y(n2777) );
AND2X1 X604 (.A(N460), .B(N154), .VDD(VDD), .VSS(VSS), .Y(n2787) );
AND2X1 X605 (.A(N443), .B(N171), .VDD(VDD), .VSS(VSS), .Y(n2797) );
AND2X1 X606 (.A(N426), .B(N188), .VDD(VDD), .VSS(VSS), .Y(n2807) );
AND2X1 X607 (.A(N409), .B(N205), .VDD(VDD), .VSS(VSS), .Y(n2817) );
AND2X1 X608 (.A(n2825), .B(n2949), .VDD(VDD), .VSS(VSS), .Y(n2827) );
AND2X1 X609 (.A(n2840), .B(n2958), .VDD(VDD), .VSS(VSS), .Y(n2950) );
AND2X1 X610 (.A(n2969), .B(n2968), .VDD(VDD), .VSS(VSS), .Y(n2962) );
AND2X1 X611 (.A(n3091), .B(n3090), .VDD(VDD), .VSS(VSS), .Y(n2957) );
AND2X1 X612 (.A(n2945), .B(n2944), .VDD(VDD), .VSS(VSS), .Y(n2973) );
AND2X1 X613 (.A(n3081), .B(n3080), .VDD(VDD), .VSS(VSS), .Y(n2972) );
AND2X1 X614 (.A(n3071), .B(n3070), .VDD(VDD), .VSS(VSS), .Y(n2974) );
AND2X1 X615 (.A(n3061), .B(n3060), .VDD(VDD), .VSS(VSS), .Y(n2976) );
AND2X1 X616 (.A(n3051), .B(n3050), .VDD(VDD), .VSS(VSS), .Y(n2978) );
AND2X1 X617 (.A(n3041), .B(n3040), .VDD(VDD), .VSS(VSS), .Y(n2980) );
AND2X1 X618 (.A(n3031), .B(n3030), .VDD(VDD), .VSS(VSS), .Y(n2982) );
AND2X1 X619 (.A(n3021), .B(n3020), .VDD(VDD), .VSS(VSS), .Y(n2984) );
AND2X1 X620 (.A(n3011), .B(n3010), .VDD(VDD), .VSS(VSS), .Y(n2986) );
AND2X1 X621 (.A(n2999), .B(n2866), .VDD(VDD), .VSS(VSS), .Y(n2867) );
AND2X1 X622 (.A(N511), .B(N86), .VDD(VDD), .VSS(VSS), .Y(n2875) );
AND2X1 X623 (.A(N494), .B(N103), .VDD(VDD), .VSS(VSS), .Y(n2885) );
AND2X1 X624 (.A(N477), .B(N120), .VDD(VDD), .VSS(VSS), .Y(n2895) );
AND2X1 X625 (.A(N460), .B(N137), .VDD(VDD), .VSS(VSS), .Y(n2905) );
AND2X1 X626 (.A(N443), .B(N154), .VDD(VDD), .VSS(VSS), .Y(n2915) );
AND2X1 X627 (.A(N426), .B(N171), .VDD(VDD), .VSS(VSS), .Y(n2925) );
AND2X1 X628 (.A(N409), .B(N188), .VDD(VDD), .VSS(VSS), .Y(n2935) );
AND2X1 X629 (.A(n2943), .B(n3079), .VDD(VDD), .VSS(VSS), .Y(n2944) );
AND2X1 X630 (.A(n2953), .B(n3089), .VDD(VDD), .VSS(VSS), .Y(n2955) );
AND2X1 X631 (.A(n2968), .B(n3098), .VDD(VDD), .VSS(VSS), .Y(n3090) );
AND2X1 X632 (.A(n3109), .B(n3108), .VDD(VDD), .VSS(VSS), .Y(n3102) );
NOR2X1 X633 (.A(n2844), .B(n2845), .Y(n2819), .VDD(VDD), .GND(VSS) );
NOR2X1 X634 (.A(n2817), .B(n2816), .Y(n2845), .VDD(VDD), .GND(VSS) );
NOR2X1 X635 (.A(n2846), .B(n2847), .Y(n2809), .VDD(VDD), .GND(VSS) );
NOR2X1 X636 (.A(n2807), .B(n2806), .Y(n2847), .VDD(VDD), .GND(VSS) );
NOR2X1 X637 (.A(n2848), .B(n2849), .Y(n2799), .VDD(VDD), .GND(VSS) );
NOR2X1 X638 (.A(n2797), .B(n2796), .Y(n2849), .VDD(VDD), .GND(VSS) );
NOR2X1 X639 (.A(n2850), .B(n2851), .Y(n2789), .VDD(VDD), .GND(VSS) );
NOR2X1 X640 (.A(n2787), .B(n2786), .Y(n2851), .VDD(VDD), .GND(VSS) );
NOR2X1 X641 (.A(n2852), .B(n2853), .Y(n2779), .VDD(VDD), .GND(VSS) );
NOR2X1 X642 (.A(n2777), .B(n2776), .Y(n2853), .VDD(VDD), .GND(VSS) );
NOR2X1 X643 (.A(n2854), .B(n2855), .Y(n2769), .VDD(VDD), .GND(VSS) );
NOR2X1 X644 (.A(n2767), .B(n2766), .Y(n2855), .VDD(VDD), .GND(VSS) );
NOR2X1 X645 (.A(n2856), .B(n2857), .Y(n2759), .VDD(VDD), .GND(VSS) );
NOR2X1 X646 (.A(n2757), .B(n2756), .Y(n2857), .VDD(VDD), .GND(VSS) );
NOR2X1 X647 (.A(n2957), .B(n2950), .Y(n2954), .VDD(VDD), .GND(VSS) );
NOR2X1 X648 (.A(n2960), .B(n2961), .Y(n2959), .VDD(VDD), .GND(VSS) );
NOR2X1 X649 (.A(n2962), .B(n2963), .Y(n2961), .VDD(VDD), .GND(VSS) );
NOR2X1 X650 (.A(N358), .B(n2843), .Y(n2960), .VDD(VDD), .GND(VSS) );
NOR2X1 X651 (.A(n2972), .B(n2973), .Y(n2947), .VDD(VDD), .GND(VSS) );
NOR2X1 X652 (.A(n2974), .B(n2975), .Y(n2937), .VDD(VDD), .GND(VSS) );
NOR2X1 X653 (.A(n2935), .B(n2934), .Y(n2975), .VDD(VDD), .GND(VSS) );
NOR2X1 X654 (.A(n2976), .B(n2977), .Y(n2927), .VDD(VDD), .GND(VSS) );
NOR2X1 X655 (.A(n2925), .B(n2924), .Y(n2977), .VDD(VDD), .GND(VSS) );
NOR2X1 X656 (.A(n2978), .B(n2979), .Y(n2917), .VDD(VDD), .GND(VSS) );
NOR2X1 X657 (.A(n2915), .B(n2914), .Y(n2979), .VDD(VDD), .GND(VSS) );
NOR2X1 X658 (.A(n2980), .B(n2981), .Y(n2907), .VDD(VDD), .GND(VSS) );
NOR2X1 X659 (.A(n2905), .B(n2904), .Y(n2981), .VDD(VDD), .GND(VSS) );
NOR2X1 X660 (.A(n2982), .B(n2983), .Y(n2897), .VDD(VDD), .GND(VSS) );
NOR2X1 X661 (.A(n2895), .B(n2894), .Y(n2983), .VDD(VDD), .GND(VSS) );
NOR2X1 X662 (.A(n2984), .B(n2985), .Y(n2887), .VDD(VDD), .GND(VSS) );
NOR2X1 X663 (.A(n2885), .B(n2884), .Y(n2985), .VDD(VDD), .GND(VSS) );
NOR2X1 X664 (.A(n2986), .B(n2987), .Y(n2877), .VDD(VDD), .GND(VSS) );
NOR2X1 X665 (.A(n2875), .B(n2874), .Y(n2987), .VDD(VDD), .GND(VSS) );
NOR2X1 X666 (.A(n3097), .B(n3090), .Y(n3094), .VDD(VDD), .GND(VSS) );
NOR2X1 X667 (.A(n3100), .B(n3101), .Y(n3099), .VDD(VDD), .GND(VSS) );
NOR2X1 X668 (.A(n3102), .B(n3103), .Y(n3101), .VDD(VDD), .GND(VSS) );
NOR2X1 X669 (.A(N341), .B(n2971), .Y(n3100), .VDD(VDD), .GND(VSS) );
NOR2X1 X670 (.A(n3112), .B(n3113), .Y(n3087), .VDD(VDD), .GND(VSS) );
NOR2X1 X671 (.A(n3085), .B(n3084), .Y(n3113), .VDD(VDD), .GND(VSS) );
NOR2X1 X672 (.A(n3114), .B(n3115), .Y(n3077), .VDD(VDD), .GND(VSS) );
NOR2X1 X673 (.A(n3075), .B(n3074), .Y(n3115), .VDD(VDD), .GND(VSS) );
NOR2X1 X674 (.A(n3116), .B(n3117), .Y(n3067), .VDD(VDD), .GND(VSS) );
NOR2X1 X675 (.A(n3065), .B(n3064), .Y(n3117), .VDD(VDD), .GND(VSS) );
NOR2X1 X676 (.A(n3118), .B(n3119), .Y(n3057), .VDD(VDD), .GND(VSS) );
NOR2X1 X677 (.A(n3055), .B(n3054), .Y(n3119), .VDD(VDD), .GND(VSS) );
NOR2X1 X678 (.A(n3120), .B(n3121), .Y(n3047), .VDD(VDD), .GND(VSS) );
NOR2X1 X679 (.A(n3045), .B(n3044), .Y(n3121), .VDD(VDD), .GND(VSS) );
NOR2X1 X680 (.A(n3122), .B(n3123), .Y(n3037), .VDD(VDD), .GND(VSS) );
NOR2X1 X681 (.A(n3035), .B(n3034), .Y(n3123), .VDD(VDD), .GND(VSS) );
NOR2X1 X682 (.A(n3124), .B(n3125), .Y(n3027), .VDD(VDD), .GND(VSS) );
NOR2X1 X683 (.A(n3025), .B(n3024), .Y(n3125), .VDD(VDD), .GND(VSS) );
NOR2X1 X684 (.A(n3126), .B(n3127), .Y(n3017), .VDD(VDD), .GND(VSS) );
NOR2X1 X685 (.A(n3015), .B(n3014), .Y(n3127), .VDD(VDD), .GND(VSS) );
NOR2X1 X686 (.A(n3128), .B(n3129), .Y(n3007), .VDD(VDD), .GND(VSS) );
NOR2X1 X687 (.A(n3005), .B(n3004), .Y(n3129), .VDD(VDD), .GND(VSS) );
NAND2X1 X688 (.A(N392), .B(N239), .Y(n2839), .VDD(VDD), .GND(VSS) );
NAND2X1 X689 (.A(N375), .B(N256), .Y(n2726), .VDD(VDD), .GND(VSS) );
NAND2X1 X690 (.A(n2840), .B(n2841), .Y(n2727), .VDD(VDD), .GND(VSS) );
NAND2X1 X691 (.A(n2842), .B(n2843), .Y(n2841), .VDD(VDD), .GND(VSS) );
NAND2X1 X692 (.A(N103), .B(N528), .Y(n2644), .VDD(VDD), .GND(VSS) );
NAND2X1 X693 (.A(n2744), .B(n2858), .Y(N6190), .VDD(VDD), .GND(VSS) );
NAND2X1 X694 (.A(n2859), .B(n2860), .Y(n2744), .VDD(VDD), .GND(VSS) );
NAND2X1 X695 (.A(n2861), .B(n2862), .Y(n2860), .VDD(VDD), .GND(VSS) );
NAND2X1 X696 (.A(n2863), .B(n2864), .Y(n2861), .VDD(VDD), .GND(VSS) );
NAND2X1 X697 (.A(n2865), .B(n2866), .Y(n2746), .VDD(VDD), .GND(VSS) );
NAND2X1 X698 (.A(n2867), .B(n2868), .Y(n2865), .VDD(VDD), .GND(VSS) );
NAND2X1 X699 (.A(n2870), .B(n2871), .Y(n2748), .VDD(VDD), .GND(VSS) );
NAND2X1 X700 (.A(n2872), .B(n2873), .Y(n2871), .VDD(VDD), .GND(VSS) );
NAND2X1 X701 (.A(n2877), .B(n2878), .Y(n2869), .VDD(VDD), .GND(VSS) );
NAND2X1 X702 (.A(n2879), .B(n2755), .Y(n2756), .VDD(VDD), .GND(VSS) );
NAND2X1 X703 (.A(n2882), .B(n2883), .Y(n2881), .VDD(VDD), .GND(VSS) );
NAND2X1 X704 (.A(n2887), .B(n2888), .Y(n2879), .VDD(VDD), .GND(VSS) );
NAND2X1 X705 (.A(n2889), .B(n2765), .Y(n2766), .VDD(VDD), .GND(VSS) );
NAND2X1 X706 (.A(n2892), .B(n2893), .Y(n2891), .VDD(VDD), .GND(VSS) );
NAND2X1 X707 (.A(n2897), .B(n2898), .Y(n2889), .VDD(VDD), .GND(VSS) );
NAND2X1 X708 (.A(n2899), .B(n2775), .Y(n2776), .VDD(VDD), .GND(VSS) );
NAND2X1 X709 (.A(n2902), .B(n2903), .Y(n2901), .VDD(VDD), .GND(VSS) );
NAND2X1 X710 (.A(n2907), .B(n2908), .Y(n2899), .VDD(VDD), .GND(VSS) );
NAND2X1 X711 (.A(n2909), .B(n2785), .Y(n2786), .VDD(VDD), .GND(VSS) );
NAND2X1 X712 (.A(n2912), .B(n2913), .Y(n2911), .VDD(VDD), .GND(VSS) );
NAND2X1 X713 (.A(n2917), .B(n2918), .Y(n2909), .VDD(VDD), .GND(VSS) );
NAND2X1 X714 (.A(n2919), .B(n2795), .Y(n2796), .VDD(VDD), .GND(VSS) );
NAND2X1 X715 (.A(n2922), .B(n2923), .Y(n2921), .VDD(VDD), .GND(VSS) );
NAND2X1 X716 (.A(n2927), .B(n2928), .Y(n2919), .VDD(VDD), .GND(VSS) );
NAND2X1 X717 (.A(n2929), .B(n2805), .Y(n2806), .VDD(VDD), .GND(VSS) );
NAND2X1 X718 (.A(n2932), .B(n2933), .Y(n2931), .VDD(VDD), .GND(VSS) );
NAND2X1 X719 (.A(n2937), .B(n2938), .Y(n2929), .VDD(VDD), .GND(VSS) );
NAND2X1 X720 (.A(n2939), .B(n2815), .Y(n2816), .VDD(VDD), .GND(VSS) );
NAND2X1 X721 (.A(n2942), .B(n2943), .Y(n2941), .VDD(VDD), .GND(VSS) );
NAND2X1 X722 (.A(n2944), .B(n2945), .Y(n2942), .VDD(VDD), .GND(VSS) );
NAND2X1 X723 (.A(n2947), .B(n2948), .Y(n2939), .VDD(VDD), .GND(VSS) );
NAND2X1 X724 (.A(N222), .B(N392), .Y(n2828), .VDD(VDD), .GND(VSS) );
NAND2X1 X725 (.A(n2952), .B(n2953), .Y(n2951), .VDD(VDD), .GND(VSS) );
NAND2X1 X726 (.A(n2954), .B(n2952), .Y(n2949), .VDD(VDD), .GND(VSS) );
NAND2X1 X727 (.A(n2955), .B(n2956), .Y(n2952), .VDD(VDD), .GND(VSS) );
NAND2X1 X728 (.A(n2959), .B(N375), .Y(n2958), .VDD(VDD), .GND(VSS) );
NAND2X1 X729 (.A(n2964), .B(n2270), .Y(n2963), .VDD(VDD), .GND(VSS) );
NAND2X1 X730 (.A(N239), .B(n2965), .Y(n2964), .VDD(VDD), .GND(VSS) );
NAND2X1 X731 (.A(n2966), .B(n2967), .Y(n2840), .VDD(VDD), .GND(VSS) );
NAND2X1 X732 (.A(N375), .B(N239), .Y(n2967), .VDD(VDD), .GND(VSS) );
NAND2X1 X733 (.A(N358), .B(N256), .Y(n2842), .VDD(VDD), .GND(VSS) );
NAND2X1 X734 (.A(n2970), .B(n2971), .Y(n2969), .VDD(VDD), .GND(VSS) );
NAND2X1 X735 (.A(N86), .B(N528), .Y(n2750), .VDD(VDD), .GND(VSS) );
NAND2X1 X736 (.A(n2862), .B(n2988), .Y(N6180), .VDD(VDD), .GND(VSS) );
NAND2X1 X737 (.A(n2989), .B(n2990), .Y(n2862), .VDD(VDD), .GND(VSS) );
NAND2X1 X738 (.A(n2991), .B(n2992), .Y(n2990), .VDD(VDD), .GND(VSS) );
NAND2X1 X739 (.A(n2993), .B(n2994), .Y(n2991), .VDD(VDD), .GND(VSS) );
NAND2X1 X740 (.A(n2995), .B(n2996), .Y(n2864), .VDD(VDD), .GND(VSS) );
NAND2X1 X741 (.A(n2997), .B(n2998), .Y(n2995), .VDD(VDD), .GND(VSS) );
NAND2X1 X742 (.A(n3000), .B(n3001), .Y(n2866), .VDD(VDD), .GND(VSS) );
NAND2X1 X743 (.A(n3002), .B(n3003), .Y(n3001), .VDD(VDD), .GND(VSS) );
NAND2X1 X744 (.A(n3007), .B(n3008), .Y(n2999), .VDD(VDD), .GND(VSS) );
NAND2X1 X745 (.A(n3009), .B(n2873), .Y(n2874), .VDD(VDD), .GND(VSS) );
NAND2X1 X746 (.A(n3012), .B(n3013), .Y(n3011), .VDD(VDD), .GND(VSS) );
NAND2X1 X747 (.A(n3017), .B(n3018), .Y(n3009), .VDD(VDD), .GND(VSS) );
NAND2X1 X748 (.A(n3019), .B(n2883), .Y(n2884), .VDD(VDD), .GND(VSS) );
NAND2X1 X749 (.A(n3022), .B(n3023), .Y(n3021), .VDD(VDD), .GND(VSS) );
NAND2X1 X750 (.A(n3027), .B(n3028), .Y(n3019), .VDD(VDD), .GND(VSS) );
NAND2X1 X751 (.A(n3029), .B(n2893), .Y(n2894), .VDD(VDD), .GND(VSS) );
NAND2X1 X752 (.A(n3032), .B(n3033), .Y(n3031), .VDD(VDD), .GND(VSS) );
NAND2X1 X753 (.A(n3037), .B(n3038), .Y(n3029), .VDD(VDD), .GND(VSS) );
NAND2X1 X754 (.A(n3039), .B(n2903), .Y(n2904), .VDD(VDD), .GND(VSS) );
NAND2X1 X755 (.A(n3042), .B(n3043), .Y(n3041), .VDD(VDD), .GND(VSS) );
NAND2X1 X756 (.A(n3047), .B(n3048), .Y(n3039), .VDD(VDD), .GND(VSS) );
NAND2X1 X757 (.A(n3049), .B(n2913), .Y(n2914), .VDD(VDD), .GND(VSS) );
NAND2X1 X758 (.A(n3052), .B(n3053), .Y(n3051), .VDD(VDD), .GND(VSS) );
NAND2X1 X759 (.A(n3057), .B(n3058), .Y(n3049), .VDD(VDD), .GND(VSS) );
NAND2X1 X760 (.A(n3059), .B(n2923), .Y(n2924), .VDD(VDD), .GND(VSS) );
NAND2X1 X761 (.A(n3062), .B(n3063), .Y(n3061), .VDD(VDD), .GND(VSS) );
NAND2X1 X762 (.A(n3067), .B(n3068), .Y(n3059), .VDD(VDD), .GND(VSS) );
NAND2X1 X763 (.A(n3069), .B(n2933), .Y(n2934), .VDD(VDD), .GND(VSS) );
NAND2X1 X764 (.A(n3072), .B(n3073), .Y(n3071), .VDD(VDD), .GND(VSS) );
NAND2X1 X765 (.A(n3077), .B(n3078), .Y(n3069), .VDD(VDD), .GND(VSS) );
NAND2X1 X766 (.A(N205), .B(N392), .Y(n2945), .VDD(VDD), .GND(VSS) );
NAND2X1 X767 (.A(n3082), .B(n3083), .Y(n3081), .VDD(VDD), .GND(VSS) );
NAND2X1 X768 (.A(n3087), .B(n3088), .Y(n3079), .VDD(VDD), .GND(VSS) );
NAND2X1 X769 (.A(N222), .B(N375), .Y(n2956), .VDD(VDD), .GND(VSS) );
NAND2X1 X770 (.A(n3092), .B(n3093), .Y(n3091), .VDD(VDD), .GND(VSS) );
NAND2X1 X771 (.A(n3094), .B(n3092), .Y(n3089), .VDD(VDD), .GND(VSS) );
NAND2X1 X772 (.A(n3095), .B(n3096), .Y(n3092), .VDD(VDD), .GND(VSS) );
NAND2X1 X773 (.A(n3099), .B(N358), .Y(n3098), .VDD(VDD), .GND(VSS) );
NAND2X1 X774 (.A(n3104), .B(n2270), .Y(n3103), .VDD(VDD), .GND(VSS) );
NAND2X1 X775 (.A(N239), .B(n3105), .Y(n3104), .VDD(VDD), .GND(VSS) );
NAND2X1 X776 (.A(n3106), .B(n3107), .Y(n2968), .VDD(VDD), .GND(VSS) );
NAND2X1 X777 (.A(N358), .B(N239), .Y(n3107), .VDD(VDD), .GND(VSS) );
NAND2X1 X778 (.A(N341), .B(N256), .Y(n2970), .VDD(VDD), .GND(VSS) );
NAND2X1 X779 (.A(n3110), .B(n3111), .Y(n3109), .VDD(VDD), .GND(VSS) );
NAND2X1 X780 (.A(N69), .B(N528), .Y(n2868), .VDD(VDD), .GND(VSS) );
NAND2X1 X781 (.A(n2992), .B(n3130), .Y(N6170), .VDD(VDD), .GND(VSS) );
NAND2X1 X782 (.A(n3131), .B(n3132), .Y(n2992), .VDD(VDD), .GND(VSS) );
NAND2X1 X783 (.A(n3133), .B(n3134), .Y(n3132), .VDD(VDD), .GND(VSS) );
NAND2X1 X784 (.A(n3135), .B(n3136), .Y(n3133), .VDD(VDD), .GND(VSS) );
NAND2X1 X785 (.A(n3137), .B(n3138), .Y(n2994), .VDD(VDD), .GND(VSS) );
INVX1 X786 (.A(n3093), .AN(n3097), .VDD(VDD), .GND(VSS) );
INVX1 X787 (.A(n3083), .AN(n3112), .VDD(VDD), .GND(VSS) );
INVX1 X788 (.A(n3073), .AN(n3114), .VDD(VDD), .GND(VSS) );
INVX1 X789 (.A(n3063), .AN(n3116), .VDD(VDD), .GND(VSS) );
INVX1 X790 (.A(n3053), .AN(n3118), .VDD(VDD), .GND(VSS) );
INVX1 X791 (.A(n3043), .AN(n3120), .VDD(VDD), .GND(VSS) );
INVX1 X792 (.A(n3033), .AN(n3122), .VDD(VDD), .GND(VSS) );
INVX1 X793 (.A(n3023), .AN(n3124), .VDD(VDD), .GND(VSS) );
INVX1 X794 (.A(n3013), .AN(n3126), .VDD(VDD), .GND(VSS) );
INVX1 X795 (.A(n3003), .AN(n3128), .VDD(VDD), .GND(VSS) );
XOR2 X796 (.A(n2998), .B(n2997), .Y(n2993), .VDD(VDD), .GND(VSS) );
XOR2 X797 (.A(n3005), .B(n3004), .Y(n3142), .VDD(VDD), .GND(VSS) );
XOR2 X798 (.A(n3004), .B(n3148), .Y(n3150), .VDD(VDD), .GND(VSS) );
XOR2 X799 (.A(n3015), .B(n3014), .Y(n3152), .VDD(VDD), .GND(VSS) );
XOR2 X800 (.A(n3014), .B(n3158), .Y(n3160), .VDD(VDD), .GND(VSS) );
XOR2 X801 (.A(n3025), .B(n3024), .Y(n3162), .VDD(VDD), .GND(VSS) );
XOR2 X802 (.A(n3024), .B(n3168), .Y(n3170), .VDD(VDD), .GND(VSS) );
XOR2 X803 (.A(n3035), .B(n3034), .Y(n3172), .VDD(VDD), .GND(VSS) );
XOR2 X804 (.A(n3034), .B(n3178), .Y(n3180), .VDD(VDD), .GND(VSS) );
XOR2 X805 (.A(n3045), .B(n3044), .Y(n3182), .VDD(VDD), .GND(VSS) );
XOR2 X806 (.A(n3044), .B(n3188), .Y(n3190), .VDD(VDD), .GND(VSS) );
XOR2 X807 (.A(n3055), .B(n3054), .Y(n3192), .VDD(VDD), .GND(VSS) );
XOR2 X808 (.A(n3054), .B(n3198), .Y(n3200), .VDD(VDD), .GND(VSS) );
XOR2 X809 (.A(n3065), .B(n3064), .Y(n3202), .VDD(VDD), .GND(VSS) );
XOR2 X810 (.A(n3064), .B(n3208), .Y(n3210), .VDD(VDD), .GND(VSS) );
XOR2 X811 (.A(n3075), .B(n3074), .Y(n3212), .VDD(VDD), .GND(VSS) );
XOR2 X812 (.A(n3074), .B(n3218), .Y(n3220), .VDD(VDD), .GND(VSS) );
XOR2 X813 (.A(n3085), .B(n3084), .Y(n3222), .VDD(VDD), .GND(VSS) );
XOR2 X814 (.A(n3084), .B(n3228), .Y(n3230), .VDD(VDD), .GND(VSS) );
XOR2 X815 (.A(n3096), .B(n3095), .Y(n3232), .VDD(VDD), .GND(VSS) );
XOR2 X816 (.A(n3238), .B(n3096), .Y(n3240), .VDD(VDD), .GND(VSS) );
XOR2 X817 (.A(n3111), .B(n3110), .Y(n3258), .VDD(VDD), .GND(VSS) );
XOR2 X818 (.A(n3135), .B(n3136), .Y(n3285), .VDD(VDD), .GND(VSS) );
XOR2 X819 (.A(n3140), .B(n3139), .Y(n3135), .VDD(VDD), .GND(VSS) );
XOR2 X820 (.A(n3147), .B(n3146), .Y(n3292), .VDD(VDD), .GND(VSS) );
XOR2 X821 (.A(n3146), .B(n3298), .Y(n3300), .VDD(VDD), .GND(VSS) );
XOR2 X822 (.A(n3157), .B(n3156), .Y(n3302), .VDD(VDD), .GND(VSS) );
XOR2 X823 (.A(n3156), .B(n3308), .Y(n3310), .VDD(VDD), .GND(VSS) );
XOR2 X824 (.A(n3167), .B(n3166), .Y(n3312), .VDD(VDD), .GND(VSS) );
XOR2 X825 (.A(n3166), .B(n3318), .Y(n3320), .VDD(VDD), .GND(VSS) );
XOR2 X826 (.A(n3177), .B(n3176), .Y(n3322), .VDD(VDD), .GND(VSS) );
XOR2 X827 (.A(n3176), .B(n3328), .Y(n3330), .VDD(VDD), .GND(VSS) );
XOR2 X828 (.A(n3187), .B(n3186), .Y(n3332), .VDD(VDD), .GND(VSS) );
XOR2 X829 (.A(n3186), .B(n3338), .Y(n3340), .VDD(VDD), .GND(VSS) );
XOR2 X830 (.A(n3197), .B(n3196), .Y(n3342), .VDD(VDD), .GND(VSS) );
XOR2 X831 (.A(n3196), .B(n3348), .Y(n3350), .VDD(VDD), .GND(VSS) );
XOR2 X832 (.A(n3207), .B(n3206), .Y(n3352), .VDD(VDD), .GND(VSS) );
XOR2 X833 (.A(n3206), .B(n3358), .Y(n3360), .VDD(VDD), .GND(VSS) );
XOR2 X834 (.A(n3217), .B(n3216), .Y(n3362), .VDD(VDD), .GND(VSS) );
XOR2 X835 (.A(n3216), .B(n3368), .Y(n3370), .VDD(VDD), .GND(VSS) );
XOR2 X836 (.A(n3227), .B(n3226), .Y(n3372), .VDD(VDD), .GND(VSS) );
XOR2 X837 (.A(n3226), .B(n3378), .Y(n3380), .VDD(VDD), .GND(VSS) );
XOR2 X838 (.A(n3237), .B(n3236), .Y(n3382), .VDD(VDD), .GND(VSS) );
XOR2 X839 (.A(n3236), .B(n3388), .Y(n3390), .VDD(VDD), .GND(VSS) );
XOR2 X840 (.A(n3248), .B(n3247), .Y(n3392), .VDD(VDD), .GND(VSS) );
XOR2 X841 (.A(n3398), .B(n3248), .Y(n3400), .VDD(VDD), .GND(VSS) );
XOR2 X842 (.A(n3263), .B(n3262), .Y(n3412), .VDD(VDD), .GND(VSS) );
OR2X1 X843 (.A(n3146), .B(n3147), .VDD(VDD), .VSS(VSS), .Y(n3144) );
OR2X1 X844 (.A(n3156), .B(n3157), .VDD(VDD), .VSS(VSS), .Y(n3154) );
OR2X1 X845 (.A(n3166), .B(n3167), .VDD(VDD), .VSS(VSS), .Y(n3164) );
OR2X1 X846 (.A(n3176), .B(n3177), .VDD(VDD), .VSS(VSS), .Y(n3174) );
OR2X1 X847 (.A(n3186), .B(n3187), .VDD(VDD), .VSS(VSS), .Y(n3184) );
OR2X1 X848 (.A(n3196), .B(n3197), .VDD(VDD), .VSS(VSS), .Y(n3194) );
OR2X1 X849 (.A(n3206), .B(n3207), .VDD(VDD), .VSS(VSS), .Y(n3204) );
OR2X1 X850 (.A(n3216), .B(n3217), .VDD(VDD), .VSS(VSS), .Y(n3214) );
OR2X1 X851 (.A(n3226), .B(n3227), .VDD(VDD), .VSS(VSS), .Y(n3224) );
OR2X1 X852 (.A(n3236), .B(n3237), .VDD(VDD), .VSS(VSS), .Y(n3234) );
OR2X1 X853 (.A(n3285), .B(n3286), .VDD(VDD), .VSS(VSS), .Y(n3284) );
OR2X1 X854 (.A(n3296), .B(n3297), .VDD(VDD), .VSS(VSS), .Y(n3294) );
OR2X1 X855 (.A(n3306), .B(n3307), .VDD(VDD), .VSS(VSS), .Y(n3304) );
OR2X1 X856 (.A(n3316), .B(n3317), .VDD(VDD), .VSS(VSS), .Y(n3314) );
OR2X1 X857 (.A(n3326), .B(n3327), .VDD(VDD), .VSS(VSS), .Y(n3324) );
OR2X1 X858 (.A(n3336), .B(n3337), .VDD(VDD), .VSS(VSS), .Y(n3334) );
OR2X1 X859 (.A(n3346), .B(n3347), .VDD(VDD), .VSS(VSS), .Y(n3344) );
OR2X1 X860 (.A(n3356), .B(n3357), .VDD(VDD), .VSS(VSS), .Y(n3354) );
OR2X1 X861 (.A(n3366), .B(n3367), .VDD(VDD), .VSS(VSS), .Y(n3364) );
OR2X1 X862 (.A(n3386), .B(n3387), .VDD(VDD), .VSS(VSS), .Y(n3384) );
OR2X1 X863 (.A(n3396), .B(n3397), .VDD(VDD), .VSS(VSS), .Y(n3394) );
OR2X1 X864 (.A(n3402), .B(n3403), .VDD(VDD), .VSS(VSS), .Y(n3245) );
AND2X1 X865 (.A(n3141), .B(n2996), .VDD(VDD), .VSS(VSS), .Y(n2997) );
AND2X1 X866 (.A(N511), .B(N69), .VDD(VDD), .VSS(VSS), .Y(n3005) );
AND2X1 X867 (.A(N494), .B(N86), .VDD(VDD), .VSS(VSS), .Y(n3015) );
AND2X1 X868 (.A(N477), .B(N103), .VDD(VDD), .VSS(VSS), .Y(n3025) );
AND2X1 X869 (.A(N460), .B(N120), .VDD(VDD), .VSS(VSS), .Y(n3035) );
AND2X1 X870 (.A(N443), .B(N137), .VDD(VDD), .VSS(VSS), .Y(n3045) );
AND2X1 X871 (.A(N426), .B(N154), .VDD(VDD), .VSS(VSS), .Y(n3055) );
AND2X1 X872 (.A(N409), .B(N171), .VDD(VDD), .VSS(VSS), .Y(n3065) );
AND2X1 X873 (.A(N392), .B(N188), .VDD(VDD), .VSS(VSS), .Y(n3075) );
AND2X1 X874 (.A(N375), .B(N205), .VDD(VDD), .VSS(VSS), .Y(n3085) );
AND2X1 X875 (.A(n3093), .B(n3241), .VDD(VDD), .VSS(VSS), .Y(n3095) );
AND2X1 X876 (.A(n3108), .B(n3250), .VDD(VDD), .VSS(VSS), .Y(n3242) );
AND2X1 X877 (.A(n3261), .B(n3260), .VDD(VDD), .VSS(VSS), .Y(n3254) );
AND2X1 X878 (.A(n3393), .B(n3392), .VDD(VDD), .VSS(VSS), .Y(n3264) );
AND2X1 X879 (.A(n3383), .B(n3382), .VDD(VDD), .VSS(VSS), .Y(n3266) );
AND2X1 X880 (.A(n3373), .B(n3372), .VDD(VDD), .VSS(VSS), .Y(n3268) );
AND2X1 X881 (.A(n3363), .B(n3362), .VDD(VDD), .VSS(VSS), .Y(n3270) );
AND2X1 X882 (.A(n3353), .B(n3352), .VDD(VDD), .VSS(VSS), .Y(n3272) );
AND2X1 X883 (.A(n3343), .B(n3342), .VDD(VDD), .VSS(VSS), .Y(n3274) );
AND2X1 X884 (.A(n3333), .B(n3332), .VDD(VDD), .VSS(VSS), .Y(n3276) );
AND2X1 X885 (.A(n3323), .B(n3322), .VDD(VDD), .VSS(VSS), .Y(n3278) );
AND2X1 X886 (.A(n3313), .B(n3312), .VDD(VDD), .VSS(VSS), .Y(n3280) );
AND2X1 X887 (.A(n3303), .B(n3302), .VDD(VDD), .VSS(VSS), .Y(n3282) );
AND2X1 X888 (.A(n3291), .B(n3138), .VDD(VDD), .VSS(VSS), .Y(n3139) );
AND2X1 X889 (.A(N511), .B(N52), .VDD(VDD), .VSS(VSS), .Y(n3147) );
AND2X1 X890 (.A(N494), .B(N69), .VDD(VDD), .VSS(VSS), .Y(n3157) );
AND2X1 X891 (.A(N477), .B(N86), .VDD(VDD), .VSS(VSS), .Y(n3167) );
AND2X1 X892 (.A(N460), .B(N103), .VDD(VDD), .VSS(VSS), .Y(n3177) );
AND2X1 X893 (.A(N443), .B(N120), .VDD(VDD), .VSS(VSS), .Y(n3187) );
AND2X1 X894 (.A(N426), .B(N137), .VDD(VDD), .VSS(VSS), .Y(n3197) );
AND2X1 X895 (.A(N409), .B(N154), .VDD(VDD), .VSS(VSS), .Y(n3207) );
AND2X1 X896 (.A(N392), .B(N171), .VDD(VDD), .VSS(VSS), .Y(n3217) );
AND2X1 X897 (.A(N375), .B(N188), .VDD(VDD), .VSS(VSS), .Y(n3227) );
AND2X1 X898 (.A(N358), .B(N205), .VDD(VDD), .VSS(VSS), .Y(n3237) );
AND2X1 X899 (.A(n3245), .B(n3401), .VDD(VDD), .VSS(VSS), .Y(n3247) );
AND2X1 X900 (.A(N290), .B(n3414), .VDD(VDD), .VSS(VSS), .Y(n3408) );
AND2X1 X901 (.A(n3415), .B(N256), .VDD(VDD), .VSS(VSS), .Y(n3414) );
AND2X1 X902 (.A(n3377), .B(n3376), .VDD(VDD), .VSS(VSS), .Y(n3424) );
NOR2X1 X903 (.A(n3249), .B(n3242), .Y(n3246), .VDD(VDD), .GND(VSS) );
NOR2X1 X904 (.A(n3252), .B(n3253), .Y(n3251), .VDD(VDD), .GND(VSS) );
NOR2X1 X905 (.A(n3254), .B(n3255), .Y(n3253), .VDD(VDD), .GND(VSS) );
NOR2X1 X906 (.A(N324), .B(n3111), .Y(n3252), .VDD(VDD), .GND(VSS) );
NOR2X1 X907 (.A(n3264), .B(n3265), .Y(n3239), .VDD(VDD), .GND(VSS) );
NOR2X1 X908 (.A(n3237), .B(n3236), .Y(n3265), .VDD(VDD), .GND(VSS) );
NOR2X1 X909 (.A(n3266), .B(n3267), .Y(n3229), .VDD(VDD), .GND(VSS) );
NOR2X1 X910 (.A(n3227), .B(n3226), .Y(n3267), .VDD(VDD), .GND(VSS) );
NOR2X1 X911 (.A(n3268), .B(n3269), .Y(n3219), .VDD(VDD), .GND(VSS) );
NOR2X1 X912 (.A(n3217), .B(n3216), .Y(n3269), .VDD(VDD), .GND(VSS) );
NOR2X1 X913 (.A(n3270), .B(n3271), .Y(n3209), .VDD(VDD), .GND(VSS) );
NOR2X1 X914 (.A(n3207), .B(n3206), .Y(n3271), .VDD(VDD), .GND(VSS) );
NOR2X1 X915 (.A(n3272), .B(n3273), .Y(n3199), .VDD(VDD), .GND(VSS) );
NOR2X1 X916 (.A(n3197), .B(n3196), .Y(n3273), .VDD(VDD), .GND(VSS) );
NOR2X1 X917 (.A(n3274), .B(n3275), .Y(n3189), .VDD(VDD), .GND(VSS) );
NOR2X1 X918 (.A(n3187), .B(n3186), .Y(n3275), .VDD(VDD), .GND(VSS) );
NOR2X1 X919 (.A(n3276), .B(n3277), .Y(n3179), .VDD(VDD), .GND(VSS) );
NOR2X1 X920 (.A(n3177), .B(n3176), .Y(n3277), .VDD(VDD), .GND(VSS) );
NOR2X1 X921 (.A(n3278), .B(n3279), .Y(n3169), .VDD(VDD), .GND(VSS) );
NOR2X1 X922 (.A(n3167), .B(n3166), .Y(n3279), .VDD(VDD), .GND(VSS) );
NOR2X1 X923 (.A(n3280), .B(n3281), .Y(n3159), .VDD(VDD), .GND(VSS) );
NOR2X1 X924 (.A(n3157), .B(n3156), .Y(n3281), .VDD(VDD), .GND(VSS) );
NOR2X1 X925 (.A(n3282), .B(n3283), .Y(n3149), .VDD(VDD), .GND(VSS) );
NOR2X1 X926 (.A(n3147), .B(n3146), .Y(n3283), .VDD(VDD), .GND(VSS) );
NOR2X1 X927 (.A(n3406), .B(n3407), .Y(n3405), .VDD(VDD), .GND(VSS) );
NOR2X1 X928 (.A(n3408), .B(n3409), .Y(n3407), .VDD(VDD), .GND(VSS) );
NOR2X1 X929 (.A(N307), .B(n3263), .Y(n3406), .VDD(VDD), .GND(VSS) );
NOR2X1 X930 (.A(n3416), .B(n3417), .Y(n3403), .VDD(VDD), .GND(VSS) );
NOR2X1 X931 (.A(n3419), .B(n3420), .Y(n3399), .VDD(VDD), .GND(VSS) );
NOR2X1 X932 (.A(n3397), .B(n3396), .Y(n3420), .VDD(VDD), .GND(VSS) );
NOR2X1 X933 (.A(n3421), .B(n3422), .Y(n3389), .VDD(VDD), .GND(VSS) );
NOR2X1 X934 (.A(n3387), .B(n3386), .Y(n3422), .VDD(VDD), .GND(VSS) );
NOR2X1 X935 (.A(n3423), .B(n3424), .Y(n3379), .VDD(VDD), .GND(VSS) );
NOR2X1 X936 (.A(n3425), .B(n3426), .Y(n3369), .VDD(VDD), .GND(VSS) );
NOR2X1 X937 (.A(n3367), .B(n3366), .Y(n3426), .VDD(VDD), .GND(VSS) );
NOR2X1 X938 (.A(n3427), .B(n3428), .Y(n3359), .VDD(VDD), .GND(VSS) );
NOR2X1 X939 (.A(n3357), .B(n3356), .Y(n3428), .VDD(VDD), .GND(VSS) );
NOR2X1 X940 (.A(n3429), .B(n3430), .Y(n3349), .VDD(VDD), .GND(VSS) );
NOR2X1 X941 (.A(n3347), .B(n3346), .Y(n3430), .VDD(VDD), .GND(VSS) );
NOR2X1 X942 (.A(n3431), .B(n3432), .Y(n3339), .VDD(VDD), .GND(VSS) );
NAND2X1 X943 (.A(n3142), .B(n3143), .Y(n2996), .VDD(VDD), .GND(VSS) );
NAND2X1 X944 (.A(n3144), .B(n3145), .Y(n3143), .VDD(VDD), .GND(VSS) );
NAND2X1 X945 (.A(n3149), .B(n3150), .Y(n3141), .VDD(VDD), .GND(VSS) );
NAND2X1 X946 (.A(n3151), .B(n3003), .Y(n3004), .VDD(VDD), .GND(VSS) );
NAND2X1 X947 (.A(n3152), .B(n3153), .Y(n3003), .VDD(VDD), .GND(VSS) );
NAND2X1 X948 (.A(n3154), .B(n3155), .Y(n3153), .VDD(VDD), .GND(VSS) );
NAND2X1 X949 (.A(n3159), .B(n3160), .Y(n3151), .VDD(VDD), .GND(VSS) );
NAND2X1 X950 (.A(n3161), .B(n3013), .Y(n3014), .VDD(VDD), .GND(VSS) );
NAND2X1 X951 (.A(n3162), .B(n3163), .Y(n3013), .VDD(VDD), .GND(VSS) );
NAND2X1 X952 (.A(n3164), .B(n3165), .Y(n3163), .VDD(VDD), .GND(VSS) );
NAND2X1 X953 (.A(n3169), .B(n3170), .Y(n3161), .VDD(VDD), .GND(VSS) );
NAND2X1 X954 (.A(n3171), .B(n3023), .Y(n3024), .VDD(VDD), .GND(VSS) );
NAND2X1 X955 (.A(n3172), .B(n3173), .Y(n3023), .VDD(VDD), .GND(VSS) );
NAND2X1 X956 (.A(n3174), .B(n3175), .Y(n3173), .VDD(VDD), .GND(VSS) );
NAND2X1 X957 (.A(n3179), .B(n3180), .Y(n3171), .VDD(VDD), .GND(VSS) );
NAND2X1 X958 (.A(n3181), .B(n3033), .Y(n3034), .VDD(VDD), .GND(VSS) );
NAND2X1 X959 (.A(n3182), .B(n3183), .Y(n3033), .VDD(VDD), .GND(VSS) );
NAND2X1 X960 (.A(n3184), .B(n3185), .Y(n3183), .VDD(VDD), .GND(VSS) );
NAND2X1 X961 (.A(n3189), .B(n3190), .Y(n3181), .VDD(VDD), .GND(VSS) );
NAND2X1 X962 (.A(n3191), .B(n3043), .Y(n3044), .VDD(VDD), .GND(VSS) );
NAND2X1 X963 (.A(n3192), .B(n3193), .Y(n3043), .VDD(VDD), .GND(VSS) );
NAND2X1 X964 (.A(n3194), .B(n3195), .Y(n3193), .VDD(VDD), .GND(VSS) );
NAND2X1 X965 (.A(n3199), .B(n3200), .Y(n3191), .VDD(VDD), .GND(VSS) );
NAND2X1 X966 (.A(n3201), .B(n3053), .Y(n3054), .VDD(VDD), .GND(VSS) );
NAND2X1 X967 (.A(n3202), .B(n3203), .Y(n3053), .VDD(VDD), .GND(VSS) );
NAND2X1 X968 (.A(n3204), .B(n3205), .Y(n3203), .VDD(VDD), .GND(VSS) );
NAND2X1 X969 (.A(n3209), .B(n3210), .Y(n3201), .VDD(VDD), .GND(VSS) );
NAND2X1 X970 (.A(n3211), .B(n3063), .Y(n3064), .VDD(VDD), .GND(VSS) );
NAND2X1 X971 (.A(n3212), .B(n3213), .Y(n3063), .VDD(VDD), .GND(VSS) );
NAND2X1 X972 (.A(n3214), .B(n3215), .Y(n3213), .VDD(VDD), .GND(VSS) );
NAND2X1 X973 (.A(n3219), .B(n3220), .Y(n3211), .VDD(VDD), .GND(VSS) );
NAND2X1 X974 (.A(n3221), .B(n3073), .Y(n3074), .VDD(VDD), .GND(VSS) );
NAND2X1 X975 (.A(n3222), .B(n3223), .Y(n3073), .VDD(VDD), .GND(VSS) );
NAND2X1 X976 (.A(n3224), .B(n3225), .Y(n3223), .VDD(VDD), .GND(VSS) );
NAND2X1 X977 (.A(n3229), .B(n3230), .Y(n3221), .VDD(VDD), .GND(VSS) );
NAND2X1 X978 (.A(n3231), .B(n3083), .Y(n3084), .VDD(VDD), .GND(VSS) );
NAND2X1 X979 (.A(n3232), .B(n3233), .Y(n3083), .VDD(VDD), .GND(VSS) );
NAND2X1 X980 (.A(n3234), .B(n3235), .Y(n3233), .VDD(VDD), .GND(VSS) );
NAND2X1 X981 (.A(n3239), .B(n3240), .Y(n3231), .VDD(VDD), .GND(VSS) );
NAND2X1 X982 (.A(N222), .B(N358), .Y(n3096), .VDD(VDD), .GND(VSS) );
NAND2X1 X983 (.A(n3242), .B(n3243), .Y(n3093), .VDD(VDD), .GND(VSS) );
NAND2X1 X984 (.A(n3244), .B(n3245), .Y(n3243), .VDD(VDD), .GND(VSS) );
NAND2X1 X985 (.A(n3246), .B(n3244), .Y(n3241), .VDD(VDD), .GND(VSS) );
NAND2X1 X986 (.A(n3247), .B(n3248), .Y(n3244), .VDD(VDD), .GND(VSS) );
NAND2X1 X987 (.A(n3251), .B(N341), .Y(n3250), .VDD(VDD), .GND(VSS) );
NAND2X1 X988 (.A(n3256), .B(n2270), .Y(n3255), .VDD(VDD), .GND(VSS) );
NAND2X1 X989 (.A(N239), .B(n3257), .Y(n3256), .VDD(VDD), .GND(VSS) );
NAND2X1 X990 (.A(n3258), .B(n3259), .Y(n3108), .VDD(VDD), .GND(VSS) );
NAND2X1 X991 (.A(N341), .B(N239), .Y(n3259), .VDD(VDD), .GND(VSS) );
NAND2X1 X992 (.A(N324), .B(N256), .Y(n3110), .VDD(VDD), .GND(VSS) );
NAND2X1 X993 (.A(n3262), .B(n3263), .Y(n3261), .VDD(VDD), .GND(VSS) );
NAND2X1 X994 (.A(N52), .B(N528), .Y(n2998), .VDD(VDD), .GND(VSS) );
NAND2X1 X995 (.A(n3134), .B(n3284), .Y(N6160), .VDD(VDD), .GND(VSS) );
NAND2X1 X996 (.A(n3285), .B(n3286), .Y(n3134), .VDD(VDD), .GND(VSS) );
NAND2X1 X997 (.A(n3287), .B(n3288), .Y(n3136), .VDD(VDD), .GND(VSS) );
NAND2X1 X998 (.A(n3289), .B(n3290), .Y(n3287), .VDD(VDD), .GND(VSS) );
NAND2X1 X999 (.A(N18), .B(N528), .Y(n3290), .VDD(VDD), .GND(VSS) );
NAND2X1 X1000 (.A(n3292), .B(n3293), .Y(n3138), .VDD(VDD), .GND(VSS) );
NAND2X1 X1001 (.A(n3294), .B(n3295), .Y(n3293), .VDD(VDD), .GND(VSS) );
NAND2X1 X1002 (.A(n3299), .B(n3300), .Y(n3291), .VDD(VDD), .GND(VSS) );
NAND2X1 X1003 (.A(n3301), .B(n3145), .Y(n3146), .VDD(VDD), .GND(VSS) );
NAND2X1 X1004 (.A(n3304), .B(n3305), .Y(n3303), .VDD(VDD), .GND(VSS) );
NAND2X1 X1005 (.A(n3309), .B(n3310), .Y(n3301), .VDD(VDD), .GND(VSS) );
NAND2X1 X1006 (.A(n3311), .B(n3155), .Y(n3156), .VDD(VDD), .GND(VSS) );
NAND2X1 X1007 (.A(n3314), .B(n3315), .Y(n3313), .VDD(VDD), .GND(VSS) );
NAND2X1 X1008 (.A(n3319), .B(n3320), .Y(n3311), .VDD(VDD), .GND(VSS) );
NAND2X1 X1009 (.A(n3321), .B(n3165), .Y(n3166), .VDD(VDD), .GND(VSS) );
NAND2X1 X1010 (.A(n3324), .B(n3325), .Y(n3323), .VDD(VDD), .GND(VSS) );
NAND2X1 X1011 (.A(n3329), .B(n3330), .Y(n3321), .VDD(VDD), .GND(VSS) );
NAND2X1 X1012 (.A(n3331), .B(n3175), .Y(n3176), .VDD(VDD), .GND(VSS) );
NAND2X1 X1013 (.A(n3334), .B(n3335), .Y(n3333), .VDD(VDD), .GND(VSS) );
NAND2X1 X1014 (.A(n3339), .B(n3340), .Y(n3331), .VDD(VDD), .GND(VSS) );
NAND2X1 X1015 (.A(n3341), .B(n3185), .Y(n3186), .VDD(VDD), .GND(VSS) );
NAND2X1 X1016 (.A(n3344), .B(n3345), .Y(n3343), .VDD(VDD), .GND(VSS) );
NAND2X1 X1017 (.A(n3349), .B(n3350), .Y(n3341), .VDD(VDD), .GND(VSS) );
NAND2X1 X1018 (.A(n3351), .B(n3195), .Y(n3196), .VDD(VDD), .GND(VSS) );
NAND2X1 X1019 (.A(n3354), .B(n3355), .Y(n3353), .VDD(VDD), .GND(VSS) );
NAND2X1 X1020 (.A(n3359), .B(n3360), .Y(n3351), .VDD(VDD), .GND(VSS) );
NAND2X1 X1021 (.A(n3361), .B(n3205), .Y(n3206), .VDD(VDD), .GND(VSS) );
NAND2X1 X1022 (.A(n3364), .B(n3365), .Y(n3363), .VDD(VDD), .GND(VSS) );
NAND2X1 X1023 (.A(n3369), .B(n3370), .Y(n3361), .VDD(VDD), .GND(VSS) );
NAND2X1 X1024 (.A(n3371), .B(n3215), .Y(n3216), .VDD(VDD), .GND(VSS) );
NAND2X1 X1025 (.A(n3374), .B(n3375), .Y(n3373), .VDD(VDD), .GND(VSS) );
NAND2X1 X1026 (.A(n3376), .B(n3377), .Y(n3374), .VDD(VDD), .GND(VSS) );
NAND2X1 X1027 (.A(n3379), .B(n3380), .Y(n3371), .VDD(VDD), .GND(VSS) );
NAND2X1 X1028 (.A(n3381), .B(n3225), .Y(n3226), .VDD(VDD), .GND(VSS) );
NAND2X1 X1029 (.A(n3384), .B(n3385), .Y(n3383), .VDD(VDD), .GND(VSS) );
NAND2X1 X1030 (.A(n3389), .B(n3390), .Y(n3381), .VDD(VDD), .GND(VSS) );
NAND2X1 X1031 (.A(n3391), .B(n3235), .Y(n3236), .VDD(VDD), .GND(VSS) );
NAND2X1 X1032 (.A(n3394), .B(n3395), .Y(n3393), .VDD(VDD), .GND(VSS) );
NAND2X1 X1033 (.A(n3399), .B(n3400), .Y(n3391), .VDD(VDD), .GND(VSS) );
NAND2X1 X1034 (.A(N222), .B(N341), .Y(n3248), .VDD(VDD), .GND(VSS) );
NAND2X1 X1035 (.A(n3403), .B(n3402), .Y(n3401), .VDD(VDD), .GND(VSS) );
NAND2X1 X1036 (.A(n3260), .B(n3404), .Y(n3402), .VDD(VDD), .GND(VSS) );
NAND2X1 X1037 (.A(n3405), .B(N324), .Y(n3404), .VDD(VDD), .GND(VSS) );
NAND2X1 X1038 (.A(n3410), .B(n2270), .Y(n3409), .VDD(VDD), .GND(VSS) );
NAND2X1 X1039 (.A(N239), .B(n3411), .Y(n3410), .VDD(VDD), .GND(VSS) );
NAND2X1 X1040 (.A(n3412), .B(n3413), .Y(n3260), .VDD(VDD), .GND(VSS) );
NAND2X1 X1041 (.A(N324), .B(N239), .Y(n3413), .VDD(VDD), .GND(VSS) );
NAND2X1 X1042 (.A(N307), .B(N256), .Y(n3262), .VDD(VDD), .GND(VSS) );
INVX1 X1043 (.A(n3418), .AN(n3417), .VDD(VDD), .GND(VSS) );
INVX1 X1044 (.A(n3395), .AN(n3419), .VDD(VDD), .GND(VSS) );
INVX1 X1045 (.A(n3385), .AN(n3421), .VDD(VDD), .GND(VSS) );
INVX1 X1046 (.A(n3375), .AN(n3423), .VDD(VDD), .GND(VSS) );
INVX1 X1047 (.A(n3365), .AN(n3425), .VDD(VDD), .GND(VSS) );
INVX1 X1048 (.A(n3355), .AN(n3427), .VDD(VDD), .GND(VSS) );
INVX1 X1049 (.A(n3345), .AN(n3429), .VDD(VDD), .GND(VSS) );
XOR2 X1050 (.A(n3445), .B(n3289), .Y(n3444), .VDD(VDD), .GND(VSS) );
XOR2 X1051 (.A(n3297), .B(n3296), .Y(n3447), .VDD(VDD), .GND(VSS) );
XOR2 X1052 (.A(n3455), .B(n3297), .Y(n3454), .VDD(VDD), .GND(VSS) );
XOR2 X1053 (.A(n3307), .B(n3306), .Y(n3458), .VDD(VDD), .GND(VSS) );
XOR2 X1054 (.A(n3306), .B(n3464), .Y(n3466), .VDD(VDD), .GND(VSS) );
XOR2 X1055 (.A(n3317), .B(n3316), .Y(n3468), .VDD(VDD), .GND(VSS) );
XOR2 X1056 (.A(n3316), .B(n3474), .Y(n3476), .VDD(VDD), .GND(VSS) );
XOR2 X1057 (.A(n3327), .B(n3326), .Y(n3478), .VDD(VDD), .GND(VSS) );
XOR2 X1058 (.A(n3326), .B(n3484), .Y(n3486), .VDD(VDD), .GND(VSS) );
XOR2 X1059 (.A(n3337), .B(n3336), .Y(n3488), .VDD(VDD), .GND(VSS) );
XOR2 X1060 (.A(n3336), .B(n3494), .Y(n3496), .VDD(VDD), .GND(VSS) );
XOR2 X1061 (.A(n3347), .B(n3346), .Y(n3498), .VDD(VDD), .GND(VSS) );
XOR2 X1062 (.A(n3346), .B(n3504), .Y(n3506), .VDD(VDD), .GND(VSS) );
XOR2 X1063 (.A(n3357), .B(n3356), .Y(n3508), .VDD(VDD), .GND(VSS) );
XOR2 X1064 (.A(n3356), .B(n3514), .Y(n3516), .VDD(VDD), .GND(VSS) );
XOR2 X1065 (.A(n3367), .B(n3366), .Y(n3518), .VDD(VDD), .GND(VSS) );
XOR2 X1066 (.A(n3366), .B(n3524), .Y(n3526), .VDD(VDD), .GND(VSS) );
XOR2 X1067 (.A(n3377), .B(n3376), .Y(n3528), .VDD(VDD), .GND(VSS) );
XOR2 X1068 (.A(n3534), .B(n3377), .Y(n3536), .VDD(VDD), .GND(VSS) );
XOR2 X1069 (.A(n3387), .B(n3386), .Y(n3538), .VDD(VDD), .GND(VSS) );
XOR2 X1070 (.A(n3386), .B(n3544), .Y(n3546), .VDD(VDD), .GND(VSS) );
XOR2 X1071 (.A(n3397), .B(n3396), .Y(n3548), .VDD(VDD), .GND(VSS) );
XOR2 X1072 (.A(n3396), .B(n3554), .Y(n3556), .VDD(VDD), .GND(VSS) );
XOR2 X1073 (.A(n3608), .B(n3607), .Y(N6123), .VDD(VDD), .GND(VSS) );
XOR2 X1074 (.A(n3452), .B(n3451), .Y(n3610), .VDD(VDD), .GND(VSS) );
XOR2 X1075 (.A(n3616), .B(n3452), .Y(n3615), .VDD(VDD), .GND(VSS) );
XOR2 X1076 (.A(n3463), .B(n3462), .Y(n3618), .VDD(VDD), .GND(VSS) );
XOR2 X1077 (.A(n3626), .B(n3463), .Y(n3625), .VDD(VDD), .GND(VSS) );
XOR2 X1078 (.A(n3473), .B(n3472), .Y(n3628), .VDD(VDD), .GND(VSS) );
XOR2 X1079 (.A(n3472), .B(n3634), .Y(n3636), .VDD(VDD), .GND(VSS) );
XOR2 X1080 (.A(n3483), .B(n3482), .Y(n3638), .VDD(VDD), .GND(VSS) );
XOR2 X1081 (.A(n3482), .B(n3644), .Y(n3646), .VDD(VDD), .GND(VSS) );
XOR2 X1082 (.A(n3493), .B(n3492), .Y(n3648), .VDD(VDD), .GND(VSS) );
XOR2 X1083 (.A(n3492), .B(n3654), .Y(n3656), .VDD(VDD), .GND(VSS) );
XOR2 X1084 (.A(n3503), .B(n3502), .Y(n3658), .VDD(VDD), .GND(VSS) );
XOR2 X1085 (.A(n3502), .B(n3664), .Y(n3666), .VDD(VDD), .GND(VSS) );
XOR2 X1086 (.A(n3513), .B(n3512), .Y(n3668), .VDD(VDD), .GND(VSS) );
XOR2 X1087 (.A(n3512), .B(n3674), .Y(n3676), .VDD(VDD), .GND(VSS) );
XOR2 X1088 (.A(n3523), .B(n3522), .Y(n3678), .VDD(VDD), .GND(VSS) );
XOR2 X1089 (.A(n3522), .B(n3684), .Y(n3686), .VDD(VDD), .GND(VSS) );
XOR2 X1090 (.A(n3533), .B(n3532), .Y(n3688), .VDD(VDD), .GND(VSS) );
XOR2 X1091 (.A(n3694), .B(n3533), .Y(n3696), .VDD(VDD), .GND(VSS) );
XOR2 X1092 (.A(n3543), .B(n3542), .Y(n3698), .VDD(VDD), .GND(VSS) );
XOR2 X1093 (.A(n3542), .B(n3704), .Y(n3706), .VDD(VDD), .GND(VSS) );
XOR2 X1094 (.A(n3553), .B(n3552), .Y(n3708), .VDD(VDD), .GND(VSS) );
XOR2 X1095 (.A(n3552), .B(n3714), .Y(n3716), .VDD(VDD), .GND(VSS) );
OR2X1 X1096 (.A(n3451), .B(n3452), .VDD(VDD), .VSS(VSS), .Y(n3449) );
OR2X1 X1097 (.A(n3462), .B(n3463), .VDD(VDD), .VSS(VSS), .Y(n3460) );
OR2X1 X1098 (.A(n3472), .B(n3473), .VDD(VDD), .VSS(VSS), .Y(n3470) );
OR2X1 X1099 (.A(n3482), .B(n3483), .VDD(VDD), .VSS(VSS), .Y(n3480) );
OR2X1 X1100 (.A(n3492), .B(n3493), .VDD(VDD), .VSS(VSS), .Y(n3490) );
OR2X1 X1101 (.A(n3502), .B(n3503), .VDD(VDD), .VSS(VSS), .Y(n3500) );
OR2X1 X1102 (.A(n3512), .B(n3513), .VDD(VDD), .VSS(VSS), .Y(n3510) );
OR2X1 X1103 (.A(n3522), .B(n3523), .VDD(VDD), .VSS(VSS), .Y(n3520) );
OR2X1 X1104 (.A(n3542), .B(n3543), .VDD(VDD), .VSS(VSS), .Y(n3540) );
OR2X1 X1105 (.A(n3552), .B(n3553), .VDD(VDD), .VSS(VSS), .Y(n3550) );
OR2X1 X1106 (.A(n3560), .B(n3561), .VDD(VDD), .VSS(VSS), .Y(n3559) );
OR2X1 X1107 (.A(n3622), .B(n3623), .VDD(VDD), .VSS(VSS), .Y(n3620) );
OR2X1 X1108 (.A(n3632), .B(n3633), .VDD(VDD), .VSS(VSS), .Y(n3630) );
OR2X1 X1109 (.A(n3642), .B(n3643), .VDD(VDD), .VSS(VSS), .Y(n3640) );
OR2X1 X1110 (.A(n3652), .B(n3653), .VDD(VDD), .VSS(VSS), .Y(n3650) );
OR2X1 X1111 (.A(n3662), .B(n3663), .VDD(VDD), .VSS(VSS), .Y(n3660) );
OR2X1 X1112 (.A(n3672), .B(n3673), .VDD(VDD), .VSS(VSS), .Y(n3670) );
OR2X1 X1113 (.A(n3682), .B(n3683), .VDD(VDD), .VSS(VSS), .Y(n3680) );
OR2X1 X1114 (.A(n3692), .B(n3693), .VDD(VDD), .VSS(VSS), .Y(n3690) );
OR2X1 X1115 (.A(n3702), .B(n3703), .VDD(VDD), .VSS(VSS), .Y(n3700) );
OR2X1 X1116 (.A(n3720), .B(n3721), .VDD(VDD), .VSS(VSS), .Y(n3719) );
AND2X1 X1117 (.A(n3499), .B(n3498), .VDD(VDD), .VSS(VSS), .Y(n3431) );
AND2X1 X1118 (.A(n3489), .B(n3488), .VDD(VDD), .VSS(VSS), .Y(n3433) );
AND2X1 X1119 (.A(n3479), .B(n3478), .VDD(VDD), .VSS(VSS), .Y(n3435) );
AND2X1 X1120 (.A(n3469), .B(n3468), .VDD(VDD), .VSS(VSS), .Y(n3437) );
AND2X1 X1121 (.A(n3459), .B(n3458), .VDD(VDD), .VSS(VSS), .Y(n3439) );
AND2X1 X1122 (.A(n3444), .B(n3443), .VDD(VDD), .VSS(VSS), .Y(n3441) );
AND2X1 X1123 (.A(n3446), .B(n3288), .VDD(VDD), .VSS(VSS), .Y(n3289) );
AND2X1 X1124 (.A(n3295), .B(n3457), .VDD(VDD), .VSS(VSS), .Y(n3455) );
AND2X1 X1125 (.A(N494), .B(N52), .VDD(VDD), .VSS(VSS), .Y(n3307) );
AND2X1 X1126 (.A(N477), .B(N69), .VDD(VDD), .VSS(VSS), .Y(n3317) );
AND2X1 X1127 (.A(N460), .B(N86), .VDD(VDD), .VSS(VSS), .Y(n3327) );
AND2X1 X1128 (.A(N443), .B(N103), .VDD(VDD), .VSS(VSS), .Y(n3337) );
AND2X1 X1129 (.A(N426), .B(N120), .VDD(VDD), .VSS(VSS), .Y(n3347) );
AND2X1 X1130 (.A(N409), .B(N137), .VDD(VDD), .VSS(VSS), .Y(n3357) );
AND2X1 X1131 (.A(N392), .B(N154), .VDD(VDD), .VSS(VSS), .Y(n3367) );
AND2X1 X1132 (.A(n3375), .B(n3537), .VDD(VDD), .VSS(VSS), .Y(n3376) );
AND2X1 X1133 (.A(N358), .B(N188), .VDD(VDD), .VSS(VSS), .Y(n3387) );
AND2X1 X1134 (.A(N341), .B(N205), .VDD(VDD), .VSS(VSS), .Y(n3397) );
AND2X1 X1135 (.A(n3418), .B(n3562), .VDD(VDD), .VSS(VSS), .Y(n3558) );
AND2X1 X1136 (.A(n3570), .B(n3569), .VDD(VDD), .VSS(VSS), .Y(n3568) );
AND2X1 X1137 (.A(n3578), .B(n3579), .VDD(VDD), .VSS(VSS), .Y(n3570) );
AND2X1 X1138 (.A(n3726), .B(n3725), .VDD(VDD), .VSS(VSS), .Y(n3560) );
AND2X1 X1139 (.A(n3719), .B(n3718), .VDD(VDD), .VSS(VSS), .Y(n3581) );
AND2X1 X1140 (.A(n3709), .B(n3708), .VDD(VDD), .VSS(VSS), .Y(n3583) );
AND2X1 X1141 (.A(n3533), .B(n3532), .VDD(VDD), .VSS(VSS), .Y(n3586) );
AND2X1 X1142 (.A(n3699), .B(n3698), .VDD(VDD), .VSS(VSS), .Y(n3585) );
AND2X1 X1143 (.A(n3689), .B(n3688), .VDD(VDD), .VSS(VSS), .Y(n3587) );
AND2X1 X1144 (.A(n3679), .B(n3678), .VDD(VDD), .VSS(VSS), .Y(n3589) );
AND2X1 X1145 (.A(n3669), .B(n3668), .VDD(VDD), .VSS(VSS), .Y(n3591) );
AND2X1 X1146 (.A(n3659), .B(n3658), .VDD(VDD), .VSS(VSS), .Y(n3593) );
AND2X1 X1147 (.A(n3649), .B(n3648), .VDD(VDD), .VSS(VSS), .Y(n3595) );
AND2X1 X1148 (.A(n3639), .B(n3638), .VDD(VDD), .VSS(VSS), .Y(n3597) );
AND2X1 X1149 (.A(n3629), .B(n3628), .VDD(VDD), .VSS(VSS), .Y(n3599) );
AND2X1 X1150 (.A(n3619), .B(n3618), .VDD(VDD), .VSS(VSS), .Y(n3601) );
AND2X1 X1151 (.A(n3604), .B(n3605), .VDD(VDD), .VSS(VSS), .Y(n3443) );
AND2X1 X1152 (.A(n3605), .B(n3609), .VDD(VDD), .VSS(VSS), .Y(n3606) );
AND2X1 X1153 (.A(n3450), .B(n3617), .VDD(VDD), .VSS(VSS), .Y(n3616) );
AND2X1 X1154 (.A(n3461), .B(n3627), .VDD(VDD), .VSS(VSS), .Y(n3626) );
AND2X1 X1155 (.A(N477), .B(N52), .VDD(VDD), .VSS(VSS), .Y(n3473) );
AND2X1 X1156 (.A(N460), .B(N69), .VDD(VDD), .VSS(VSS), .Y(n3483) );
AND2X1 X1157 (.A(N443), .B(N86), .VDD(VDD), .VSS(VSS), .Y(n3493) );
AND2X1 X1158 (.A(N426), .B(N103), .VDD(VDD), .VSS(VSS), .Y(n3503) );
AND2X1 X1159 (.A(N409), .B(N120), .VDD(VDD), .VSS(VSS), .Y(n3513) );
AND2X1 X1160 (.A(N392), .B(N137), .VDD(VDD), .VSS(VSS), .Y(n3523) );
AND2X1 X1161 (.A(n3531), .B(n3697), .VDD(VDD), .VSS(VSS), .Y(n3532) );
AND2X1 X1162 (.A(N358), .B(N171), .VDD(VDD), .VSS(VSS), .Y(n3543) );
AND2X1 X1163 (.A(N341), .B(N188), .VDD(VDD), .VSS(VSS), .Y(n3553) );
AND2X1 X1164 (.A(n3580), .B(n3722), .VDD(VDD), .VSS(VSS), .Y(n3718) );
NOR2X1 X1165 (.A(n3337), .B(n3336), .Y(n3432), .VDD(VDD), .GND(VSS) );
NOR2X1 X1166 (.A(n3433), .B(n3434), .Y(n3329), .VDD(VDD), .GND(VSS) );
NOR2X1 X1167 (.A(n3327), .B(n3326), .Y(n3434), .VDD(VDD), .GND(VSS) );
NOR2X1 X1168 (.A(n3435), .B(n3436), .Y(n3319), .VDD(VDD), .GND(VSS) );
NOR2X1 X1169 (.A(n3317), .B(n3316), .Y(n3436), .VDD(VDD), .GND(VSS) );
NOR2X1 X1170 (.A(n3437), .B(n3438), .Y(n3309), .VDD(VDD), .GND(VSS) );
NOR2X1 X1171 (.A(n3307), .B(n3306), .Y(n3438), .VDD(VDD), .GND(VSS) );
NOR2X1 X1172 (.A(n3439), .B(n3440), .Y(n3299), .VDD(VDD), .GND(VSS) );
NOR2X1 X1173 (.A(n3297), .B(n3296), .Y(n3440), .VDD(VDD), .GND(VSS) );
NOR2X1 X1174 (.A(n3441), .B(n3442), .Y(N6150), .VDD(VDD), .GND(VSS) );
NOR2X1 X1175 (.A(n3443), .B(n3444), .Y(n3442), .VDD(VDD), .GND(VSS) );
NOR2X1 X1176 (.A(n3456), .B(n2232), .Y(n3297), .VDD(VDD), .GND(VSS) );
NOR2X1 X1177 (.A(n3565), .B(n3257), .Y(n3567), .VDD(VDD), .GND(VSS) );
NOR2X1 X1178 (.A(n3568), .B(n3416), .Y(n3565), .VDD(VDD), .GND(VSS) );
NOR2X1 X1179 (.A(n3569), .B(n3570), .Y(n3416), .VDD(VDD), .GND(VSS) );
NOR2X1 X1180 (.A(n3577), .B(n2275), .Y(n3575), .VDD(VDD), .GND(VSS) );
NOR2X1 X1181 (.A(n2228), .B(n3411), .Y(n3577), .VDD(VDD), .GND(VSS) );
NOR2X1 X1182 (.A(n3561), .B(n3560), .Y(n3563), .VDD(VDD), .GND(VSS) );
NOR2X1 X1183 (.A(n3581), .B(n3582), .Y(n3555), .VDD(VDD), .GND(VSS) );
NOR2X1 X1184 (.A(n3553), .B(n3552), .Y(n3582), .VDD(VDD), .GND(VSS) );
NOR2X1 X1185 (.A(n3583), .B(n3584), .Y(n3545), .VDD(VDD), .GND(VSS) );
NOR2X1 X1186 (.A(n3543), .B(n3542), .Y(n3584), .VDD(VDD), .GND(VSS) );
NOR2X1 X1187 (.A(n3585), .B(n3586), .Y(n3535), .VDD(VDD), .GND(VSS) );
NOR2X1 X1188 (.A(n3587), .B(n3588), .Y(n3525), .VDD(VDD), .GND(VSS) );
NOR2X1 X1189 (.A(n3523), .B(n3522), .Y(n3588), .VDD(VDD), .GND(VSS) );
NOR2X1 X1190 (.A(n3589), .B(n3590), .Y(n3515), .VDD(VDD), .GND(VSS) );
NOR2X1 X1191 (.A(n3513), .B(n3512), .Y(n3590), .VDD(VDD), .GND(VSS) );
NOR2X1 X1192 (.A(n3591), .B(n3592), .Y(n3505), .VDD(VDD), .GND(VSS) );
NOR2X1 X1193 (.A(n3503), .B(n3502), .Y(n3592), .VDD(VDD), .GND(VSS) );
NOR2X1 X1194 (.A(n3593), .B(n3594), .Y(n3495), .VDD(VDD), .GND(VSS) );
NOR2X1 X1195 (.A(n3493), .B(n3492), .Y(n3594), .VDD(VDD), .GND(VSS) );
NOR2X1 X1196 (.A(n3595), .B(n3596), .Y(n3485), .VDD(VDD), .GND(VSS) );
NOR2X1 X1197 (.A(n3483), .B(n3482), .Y(n3596), .VDD(VDD), .GND(VSS) );
NOR2X1 X1198 (.A(n3597), .B(n3598), .Y(n3475), .VDD(VDD), .GND(VSS) );
NOR2X1 X1199 (.A(n3473), .B(n3472), .Y(n3598), .VDD(VDD), .GND(VSS) );
NOR2X1 X1200 (.A(n3599), .B(n3600), .Y(n3465), .VDD(VDD), .GND(VSS) );
NOR2X1 X1201 (.A(n3463), .B(n3462), .Y(n3600), .VDD(VDD), .GND(VSS) );
NOR2X1 X1202 (.A(n3601), .B(n3602), .Y(n3453), .VDD(VDD), .GND(VSS) );
NOR2X1 X1203 (.A(n3452), .B(n3451), .Y(n3602), .VDD(VDD), .GND(VSS) );
NOR2X1 X1204 (.A(n3603), .B(n2205), .Y(n3445), .VDD(VDD), .GND(VSS) );
NOR2X1 X1205 (.A(n3603), .B(n2232), .Y(n3452), .VDD(VDD), .GND(VSS) );
NOR2X1 X1206 (.A(n3456), .B(n2271), .Y(n3463), .VDD(VDD), .GND(VSS) );
NAND2X1 X1207 (.A(N35), .B(N528), .Y(n3140), .VDD(VDD), .GND(VSS) );
NAND2X1 X1208 (.A(n3447), .B(n3448), .Y(n3288), .VDD(VDD), .GND(VSS) );
NAND2X1 X1209 (.A(n3449), .B(n3450), .Y(n3448), .VDD(VDD), .GND(VSS) );
NAND2X1 X1210 (.A(n3453), .B(n3454), .Y(n3446), .VDD(VDD), .GND(VSS) );
NAND2X1 X1211 (.A(n3460), .B(n3461), .Y(n3459), .VDD(VDD), .GND(VSS) );
NAND2X1 X1212 (.A(n3465), .B(n3466), .Y(n3457), .VDD(VDD), .GND(VSS) );
NAND2X1 X1213 (.A(n3467), .B(n3305), .Y(n3306), .VDD(VDD), .GND(VSS) );
NAND2X1 X1214 (.A(n3470), .B(n3471), .Y(n3469), .VDD(VDD), .GND(VSS) );
NAND2X1 X1215 (.A(n3475), .B(n3476), .Y(n3467), .VDD(VDD), .GND(VSS) );
NAND2X1 X1216 (.A(n3477), .B(n3315), .Y(n3316), .VDD(VDD), .GND(VSS) );
NAND2X1 X1217 (.A(n3480), .B(n3481), .Y(n3479), .VDD(VDD), .GND(VSS) );
NAND2X1 X1218 (.A(n3485), .B(n3486), .Y(n3477), .VDD(VDD), .GND(VSS) );
NAND2X1 X1219 (.A(n3487), .B(n3325), .Y(n3326), .VDD(VDD), .GND(VSS) );
NAND2X1 X1220 (.A(n3490), .B(n3491), .Y(n3489), .VDD(VDD), .GND(VSS) );
NAND2X1 X1221 (.A(n3495), .B(n3496), .Y(n3487), .VDD(VDD), .GND(VSS) );
NAND2X1 X1222 (.A(n3497), .B(n3335), .Y(n3336), .VDD(VDD), .GND(VSS) );
NAND2X1 X1223 (.A(n3500), .B(n3501), .Y(n3499), .VDD(VDD), .GND(VSS) );
NAND2X1 X1224 (.A(n3505), .B(n3506), .Y(n3497), .VDD(VDD), .GND(VSS) );
NAND2X1 X1225 (.A(n3507), .B(n3345), .Y(n3346), .VDD(VDD), .GND(VSS) );
NAND2X1 X1226 (.A(n3508), .B(n3509), .Y(n3345), .VDD(VDD), .GND(VSS) );
NAND2X1 X1227 (.A(n3510), .B(n3511), .Y(n3509), .VDD(VDD), .GND(VSS) );
NAND2X1 X1228 (.A(n3515), .B(n3516), .Y(n3507), .VDD(VDD), .GND(VSS) );
NAND2X1 X1229 (.A(n3517), .B(n3355), .Y(n3356), .VDD(VDD), .GND(VSS) );
NAND2X1 X1230 (.A(n3518), .B(n3519), .Y(n3355), .VDD(VDD), .GND(VSS) );
NAND2X1 X1231 (.A(n3520), .B(n3521), .Y(n3519), .VDD(VDD), .GND(VSS) );
NAND2X1 X1232 (.A(n3525), .B(n3526), .Y(n3517), .VDD(VDD), .GND(VSS) );
NAND2X1 X1233 (.A(n3527), .B(n3365), .Y(n3366), .VDD(VDD), .GND(VSS) );
NAND2X1 X1234 (.A(n3528), .B(n3529), .Y(n3365), .VDD(VDD), .GND(VSS) );
NAND2X1 X1235 (.A(n3530), .B(n3531), .Y(n3529), .VDD(VDD), .GND(VSS) );
NAND2X1 X1236 (.A(n3532), .B(n3533), .Y(n3530), .VDD(VDD), .GND(VSS) );
NAND2X1 X1237 (.A(n3535), .B(n3536), .Y(n3527), .VDD(VDD), .GND(VSS) );
NAND2X1 X1238 (.A(N171), .B(N375), .Y(n3377), .VDD(VDD), .GND(VSS) );
NAND2X1 X1239 (.A(n3538), .B(n3539), .Y(n3375), .VDD(VDD), .GND(VSS) );
NAND2X1 X1240 (.A(n3540), .B(n3541), .Y(n3539), .VDD(VDD), .GND(VSS) );
NAND2X1 X1241 (.A(n3545), .B(n3546), .Y(n3537), .VDD(VDD), .GND(VSS) );
NAND2X1 X1242 (.A(n3547), .B(n3385), .Y(n3386), .VDD(VDD), .GND(VSS) );
NAND2X1 X1243 (.A(n3548), .B(n3549), .Y(n3385), .VDD(VDD), .GND(VSS) );
NAND2X1 X1244 (.A(n3550), .B(n3551), .Y(n3549), .VDD(VDD), .GND(VSS) );
NAND2X1 X1245 (.A(n3555), .B(n3556), .Y(n3547), .VDD(VDD), .GND(VSS) );
NAND2X1 X1246 (.A(n3557), .B(n3395), .Y(n3396), .VDD(VDD), .GND(VSS) );
NAND2X1 X1247 (.A(n3558), .B(n3559), .Y(n3395), .VDD(VDD), .GND(VSS) );
NAND2X1 X1248 (.A(n3563), .B(n3564), .Y(n3557), .VDD(VDD), .GND(VSS) );
NAND2X1 X1249 (.A(n3562), .B(n3418), .Y(n3564), .VDD(VDD), .GND(VSS) );
NAND2X1 X1250 (.A(n3565), .B(n3566), .Y(n3418), .VDD(VDD), .GND(VSS) );
NAND2X1 X1251 (.A(N222), .B(N324), .Y(n3566), .VDD(VDD), .GND(VSS) );
NAND2X1 X1252 (.A(n3567), .B(N222), .Y(n3562), .VDD(VDD), .GND(VSS) );
NAND2X1 X1253 (.A(n3415), .B(n3571), .Y(n3569), .VDD(VDD), .GND(VSS) );
NAND2X1 X1254 (.A(N307), .B(n3572), .Y(n3571), .VDD(VDD), .GND(VSS) );
NAND2X1 X1255 (.A(n2270), .B(n3573), .Y(n3572), .VDD(VDD), .GND(VSS) );
NAND2X1 X1256 (.A(N239), .B(n3574), .Y(n3573), .VDD(VDD), .GND(VSS) );
NAND2X1 X1257 (.A(N239), .B(n2275), .Y(n2270), .VDD(VDD), .GND(VSS) );
NAND2X1 X1258 (.A(n3575), .B(n3576), .Y(n3415), .VDD(VDD), .GND(VSS) );
NAND2X1 X1259 (.A(n3606), .B(n3607), .Y(n3604), .VDD(VDD), .GND(VSS) );
NAND2X1 X1260 (.A(N1), .B(N528), .Y(n3607), .VDD(VDD), .GND(VSS) );
NAND2X1 X1261 (.A(n3610), .B(n3611), .Y(n3605), .VDD(VDD), .GND(VSS) );
NAND2X1 X1262 (.A(n3612), .B(n3613), .Y(n3611), .VDD(VDD), .GND(VSS) );
NAND2X1 X1263 (.A(n3614), .B(n3615), .Y(n3609), .VDD(VDD), .GND(VSS) );
NAND2X1 X1264 (.A(n3620), .B(n3621), .Y(n3619), .VDD(VDD), .GND(VSS) );
NAND2X1 X1265 (.A(n3624), .B(n3625), .Y(n3617), .VDD(VDD), .GND(VSS) );
NAND2X1 X1266 (.A(n3630), .B(n3631), .Y(n3629), .VDD(VDD), .GND(VSS) );
NAND2X1 X1267 (.A(n3635), .B(n3636), .Y(n3627), .VDD(VDD), .GND(VSS) );
NAND2X1 X1268 (.A(n3637), .B(n3471), .Y(n3472), .VDD(VDD), .GND(VSS) );
NAND2X1 X1269 (.A(n3640), .B(n3641), .Y(n3639), .VDD(VDD), .GND(VSS) );
NAND2X1 X1270 (.A(n3645), .B(n3646), .Y(n3637), .VDD(VDD), .GND(VSS) );
NAND2X1 X1271 (.A(n3647), .B(n3481), .Y(n3482), .VDD(VDD), .GND(VSS) );
NAND2X1 X1272 (.A(n3650), .B(n3651), .Y(n3649), .VDD(VDD), .GND(VSS) );
NAND2X1 X1273 (.A(n3655), .B(n3656), .Y(n3647), .VDD(VDD), .GND(VSS) );
NAND2X1 X1274 (.A(n3657), .B(n3491), .Y(n3492), .VDD(VDD), .GND(VSS) );
NAND2X1 X1275 (.A(n3660), .B(n3661), .Y(n3659), .VDD(VDD), .GND(VSS) );
NAND2X1 X1276 (.A(n3665), .B(n3666), .Y(n3657), .VDD(VDD), .GND(VSS) );
NAND2X1 X1277 (.A(n3667), .B(n3501), .Y(n3502), .VDD(VDD), .GND(VSS) );
NAND2X1 X1278 (.A(n3670), .B(n3671), .Y(n3669), .VDD(VDD), .GND(VSS) );
NAND2X1 X1279 (.A(n3675), .B(n3676), .Y(n3667), .VDD(VDD), .GND(VSS) );
NAND2X1 X1280 (.A(n3677), .B(n3511), .Y(n3512), .VDD(VDD), .GND(VSS) );
NAND2X1 X1281 (.A(n3680), .B(n3681), .Y(n3679), .VDD(VDD), .GND(VSS) );
NAND2X1 X1282 (.A(n3685), .B(n3686), .Y(n3677), .VDD(VDD), .GND(VSS) );
NAND2X1 X1283 (.A(n3687), .B(n3521), .Y(n3522), .VDD(VDD), .GND(VSS) );
NAND2X1 X1284 (.A(n3690), .B(n3691), .Y(n3689), .VDD(VDD), .GND(VSS) );
NAND2X1 X1285 (.A(n3695), .B(n3696), .Y(n3687), .VDD(VDD), .GND(VSS) );
NAND2X1 X1286 (.A(N154), .B(N375), .Y(n3533), .VDD(VDD), .GND(VSS) );
NAND2X1 X1287 (.A(n3700), .B(n3701), .Y(n3699), .VDD(VDD), .GND(VSS) );
NAND2X1 X1288 (.A(n3705), .B(n3706), .Y(n3697), .VDD(VDD), .GND(VSS) );
NAND2X1 X1289 (.A(n3707), .B(n3541), .Y(n3542), .VDD(VDD), .GND(VSS) );
NAND2X1 X1290 (.A(n3710), .B(n3711), .Y(n3709), .VDD(VDD), .GND(VSS) );
NAND2X1 X1291 (.A(n3712), .B(n3713), .Y(n3710), .VDD(VDD), .GND(VSS) );
NAND2X1 X1292 (.A(n3715), .B(n3716), .Y(n3707), .VDD(VDD), .GND(VSS) );
NAND2X1 X1293 (.A(n3717), .B(n3551), .Y(n3552), .VDD(VDD), .GND(VSS) );
NAND2X1 X1294 (.A(n3723), .B(n3724), .Y(n3717), .VDD(VDD), .GND(VSS) );
NAND2X1 X1295 (.A(n3722), .B(n3580), .Y(n3724), .VDD(VDD), .GND(VSS) );
NAND2X1 X1296 (.A(N205), .B(N324), .Y(n3726), .VDD(VDD), .GND(VSS) );
NAND2X1 X1297 (.A(n3727), .B(N205), .Y(n3722), .VDD(VDD), .GND(VSS) );
INVX1 X1298 (.A(N528), .AN(n2205), .VDD(VDD), .GND(VSS) );
XOR2 X1299 (.A(n3623), .B(n3622), .Y(n3775), .VDD(VDD), .GND(VSS) );
XOR2 X1300 (.A(n3783), .B(n3623), .Y(n3782), .VDD(VDD), .GND(VSS) );
XOR2 X1301 (.A(n3633), .B(n3632), .Y(n3785), .VDD(VDD), .GND(VSS) );
XOR2 X1302 (.A(n3793), .B(n3633), .Y(n3792), .VDD(VDD), .GND(VSS) );
XOR2 X1303 (.A(n3643), .B(n3642), .Y(n3795), .VDD(VDD), .GND(VSS) );
XOR2 X1304 (.A(n3642), .B(n3801), .Y(n3803), .VDD(VDD), .GND(VSS) );
XOR2 X1305 (.A(n3653), .B(n3652), .Y(n3805), .VDD(VDD), .GND(VSS) );
XOR2 X1306 (.A(n3652), .B(n3811), .Y(n3813), .VDD(VDD), .GND(VSS) );
XOR2 X1307 (.A(n3663), .B(n3662), .Y(n3815), .VDD(VDD), .GND(VSS) );
XOR2 X1308 (.A(n3662), .B(n3821), .Y(n3823), .VDD(VDD), .GND(VSS) );
XOR2 X1309 (.A(n3673), .B(n3672), .Y(n3825), .VDD(VDD), .GND(VSS) );
XOR2 X1310 (.A(n3672), .B(n3831), .Y(n3833), .VDD(VDD), .GND(VSS) );
XOR2 X1311 (.A(n3683), .B(n3682), .Y(n3835), .VDD(VDD), .GND(VSS) );
XOR2 X1312 (.A(n3682), .B(n3841), .Y(n3843), .VDD(VDD), .GND(VSS) );
XOR2 X1313 (.A(n3693), .B(n3692), .Y(n3845), .VDD(VDD), .GND(VSS) );
XOR2 X1314 (.A(n3692), .B(n3851), .Y(n3853), .VDD(VDD), .GND(VSS) );
XOR2 X1315 (.A(n3703), .B(n3702), .Y(n3855), .VDD(VDD), .GND(VSS) );
XOR2 X1316 (.A(n3702), .B(n3861), .Y(n3863), .VDD(VDD), .GND(VSS) );
XOR2 X1317 (.A(n3713), .B(n3712), .Y(n3865), .VDD(VDD), .GND(VSS) );
XOR2 X1318 (.A(n3871), .B(n3713), .Y(n3873), .VDD(VDD), .GND(VSS) );
XOR2 X1319 (.A(n3928), .B(n3780), .Y(N5672), .VDD(VDD), .GND(VSS) );
XOR2 X1320 (.A(n3790), .B(n3789), .Y(n3931), .VDD(VDD), .GND(VSS) );
XOR2 X1321 (.A(n3925), .B(n3790), .Y(n3938), .VDD(VDD), .GND(VSS) );
XOR2 X1322 (.A(n3800), .B(n3799), .Y(n3940), .VDD(VDD), .GND(VSS) );
XOR2 X1323 (.A(n3921), .B(n3800), .Y(n3947), .VDD(VDD), .GND(VSS) );
XOR2 X1324 (.A(n3810), .B(n3809), .Y(n3949), .VDD(VDD), .GND(VSS) );
XOR2 X1325 (.A(n3955), .B(n3810), .Y(n3957), .VDD(VDD), .GND(VSS) );
XOR2 X1326 (.A(n3820), .B(n3819), .Y(n3959), .VDD(VDD), .GND(VSS) );
XOR2 X1327 (.A(n3965), .B(n3820), .Y(n3967), .VDD(VDD), .GND(VSS) );
XOR2 X1328 (.A(n3830), .B(n3829), .Y(n3969), .VDD(VDD), .GND(VSS) );
XOR2 X1329 (.A(n3975), .B(n3830), .Y(n3977), .VDD(VDD), .GND(VSS) );
XOR2 X1330 (.A(n3840), .B(n3839), .Y(n3979), .VDD(VDD), .GND(VSS) );
XOR2 X1331 (.A(n3985), .B(n3840), .Y(n3987), .VDD(VDD), .GND(VSS) );
XOR2 X1332 (.A(n3850), .B(n3849), .Y(n3989), .VDD(VDD), .GND(VSS) );
XOR2 X1333 (.A(n3995), .B(n3850), .Y(n3997), .VDD(VDD), .GND(VSS) );
XOR2 X1334 (.A(n3860), .B(n3859), .Y(n3999), .VDD(VDD), .GND(VSS) );
XOR2 X1335 (.A(n3859), .B(n4005), .Y(n4007), .VDD(VDD), .GND(VSS) );
XOR2 X1336 (.A(n3870), .B(n3869), .Y(n4009), .VDD(VDD), .GND(VSS) );
XOR2 X1337 (.A(n4015), .B(n3870), .Y(n4017), .VDD(VDD), .GND(VSS) );
OR2X1 X1338 (.A(n3779), .B(n3780), .VDD(VDD), .VSS(VSS), .Y(n3777) );
OR2X1 X1339 (.A(n3859), .B(n3860), .VDD(VDD), .VSS(VSS), .Y(n3857) );
OR2X1 X1340 (.A(n3877), .B(n3878), .VDD(VDD), .VSS(VSS), .Y(n3876) );
OR2X1 X1341 (.A(n3893), .B(n3736), .VDD(VDD), .VSS(VSS), .Y(n3892) );
OR2X1 X1342 (.A(n3935), .B(n3936), .VDD(VDD), .VSS(VSS), .Y(n3933) );
OR2X1 X1343 (.A(n4003), .B(n4004), .VDD(VDD), .VSS(VSS), .Y(n4001) );
OR2X1 X1344 (.A(n4021), .B(n4022), .VDD(VDD), .VSS(VSS), .Y(n4020) );
AND2X1 X1345 (.A(n3730), .B(n3729), .VDD(VDD), .VSS(VSS), .Y(n3728) );
AND2X1 X1346 (.A(n3579), .B(n3735), .VDD(VDD), .VSS(VSS), .Y(n3733) );
AND2X1 X1347 (.A(n3737), .B(N290), .VDD(VDD), .VSS(VSS), .Y(n3576) );
AND2X1 X1348 (.A(n3747), .B(n3748), .VDD(VDD), .VSS(VSS), .Y(n3730) );
AND2X1 X1349 (.A(n3883), .B(n3882), .VDD(VDD), .VSS(VSS), .Y(n3720) );
AND2X1 X1350 (.A(n3713), .B(n3712), .VDD(VDD), .VSS(VSS), .Y(n3751) );
AND2X1 X1351 (.A(n3876), .B(n3875), .VDD(VDD), .VSS(VSS), .Y(n3750) );
AND2X1 X1352 (.A(n3866), .B(n3865), .VDD(VDD), .VSS(VSS), .Y(n3752) );
AND2X1 X1353 (.A(n3856), .B(n3855), .VDD(VDD), .VSS(VSS), .Y(n3754) );
AND2X1 X1354 (.A(n3846), .B(n3845), .VDD(VDD), .VSS(VSS), .Y(n3756) );
AND2X1 X1355 (.A(n3836), .B(n3835), .VDD(VDD), .VSS(VSS), .Y(n3758) );
AND2X1 X1356 (.A(n3826), .B(n3825), .VDD(VDD), .VSS(VSS), .Y(n3760) );
AND2X1 X1357 (.A(n3816), .B(n3815), .VDD(VDD), .VSS(VSS), .Y(n3762) );
AND2X1 X1358 (.A(n3806), .B(n3805), .VDD(VDD), .VSS(VSS), .Y(n3764) );
AND2X1 X1359 (.A(n3796), .B(n3795), .VDD(VDD), .VSS(VSS), .Y(n3766) );
AND2X1 X1360 (.A(n3786), .B(n3785), .VDD(VDD), .VSS(VSS), .Y(n3768) );
AND2X1 X1361 (.A(n3613), .B(n3612), .VDD(VDD), .VSS(VSS), .Y(n3614) );
AND2X1 X1362 (.A(n3774), .B(n3613), .VDD(VDD), .VSS(VSS), .Y(n3772) );
AND2X1 X1363 (.A(n3621), .B(n3784), .VDD(VDD), .VSS(VSS), .Y(n3783) );
AND2X1 X1364 (.A(n3631), .B(n3794), .VDD(VDD), .VSS(VSS), .Y(n3793) );
AND2X1 X1365 (.A(N460), .B(N52), .VDD(VDD), .VSS(VSS), .Y(n3643) );
AND2X1 X1366 (.A(N443), .B(N69), .VDD(VDD), .VSS(VSS), .Y(n3653) );
AND2X1 X1367 (.A(N426), .B(N86), .VDD(VDD), .VSS(VSS), .Y(n3663) );
AND2X1 X1368 (.A(N409), .B(N103), .VDD(VDD), .VSS(VSS), .Y(n3673) );
AND2X1 X1369 (.A(N392), .B(N120), .VDD(VDD), .VSS(VSS), .Y(n3683) );
AND2X1 X1370 (.A(N375), .B(N137), .VDD(VDD), .VSS(VSS), .Y(n3693) );
AND2X1 X1371 (.A(N358), .B(N154), .VDD(VDD), .VSS(VSS), .Y(n3703) );
AND2X1 X1372 (.A(n3711), .B(n3874), .VDD(VDD), .VSS(VSS), .Y(n3712) );
AND2X1 X1373 (.A(n3749), .B(n3879), .VDD(VDD), .VSS(VSS), .Y(n3875) );
AND2X1 X1374 (.A(n3887), .B(n3886), .VDD(VDD), .VSS(VSS), .Y(n3885) );
AND2X1 X1375 (.A(n3748), .B(n3892), .VDD(VDD), .VSS(VSS), .Y(n3890) );
AND2X1 X1376 (.A(N222), .B(n3897), .VDD(VDD), .VSS(VSS), .Y(n3736) );
AND2X1 X1377 (.A(n3901), .B(n3902), .VDD(VDD), .VSS(VSS), .Y(n3887) );
AND2X1 X1378 (.A(n4027), .B(n4026), .VDD(VDD), .VSS(VSS), .Y(n3877) );
AND2X1 X1379 (.A(n3870), .B(n3869), .VDD(VDD), .VSS(VSS), .Y(n3905) );
AND2X1 X1380 (.A(n4020), .B(n4019), .VDD(VDD), .VSS(VSS), .Y(n3904) );
AND2X1 X1381 (.A(n4010), .B(n4009), .VDD(VDD), .VSS(VSS), .Y(n3906) );
AND2X1 X1382 (.A(n3850), .B(n3849), .VDD(VDD), .VSS(VSS), .Y(n3909) );
AND2X1 X1383 (.A(n4000), .B(n3999), .VDD(VDD), .VSS(VSS), .Y(n3908) );
AND2X1 X1384 (.A(n3840), .B(n3839), .VDD(VDD), .VSS(VSS), .Y(n3911) );
AND2X1 X1385 (.A(n3990), .B(n3989), .VDD(VDD), .VSS(VSS), .Y(n3910) );
AND2X1 X1386 (.A(n3830), .B(n3829), .VDD(VDD), .VSS(VSS), .Y(n3913) );
AND2X1 X1387 (.A(n3980), .B(n3979), .VDD(VDD), .VSS(VSS), .Y(n3912) );
AND2X1 X1388 (.A(n3820), .B(n3819), .VDD(VDD), .VSS(VSS), .Y(n3915) );
AND2X1 X1389 (.A(n3970), .B(n3969), .VDD(VDD), .VSS(VSS), .Y(n3914) );
AND2X1 X1390 (.A(n3810), .B(n3809), .VDD(VDD), .VSS(VSS), .Y(n3917) );
AND2X1 X1391 (.A(n3960), .B(n3959), .VDD(VDD), .VSS(VSS), .Y(n3916) );
AND2X1 X1392 (.A(N460), .B(N35), .VDD(VDD), .VSS(VSS), .Y(n3920) );
AND2X1 X1393 (.A(n3950), .B(n3949), .VDD(VDD), .VSS(VSS), .Y(n3918) );
AND2X1 X1394 (.A(N477), .B(N18), .VDD(VDD), .VSS(VSS), .Y(n3924) );
AND2X1 X1395 (.A(n3941), .B(n3940), .VDD(VDD), .VSS(VSS), .Y(n3922) );
AND2X1 X1396 (.A(n3932), .B(n3931), .VDD(VDD), .VSS(VSS), .Y(n3926) );
AND2X1 X1397 (.A(n3778), .B(n3930), .VDD(VDD), .VSS(VSS), .Y(n3928) );
AND2X1 X1398 (.A(n3788), .B(n3939), .VDD(VDD), .VSS(VSS), .Y(n3789) );
AND2X1 X1399 (.A(n3798), .B(n3948), .VDD(VDD), .VSS(VSS), .Y(n3799) );
AND2X1 X1400 (.A(n3808), .B(n3958), .VDD(VDD), .VSS(VSS), .Y(n3809) );
AND2X1 X1401 (.A(n3818), .B(n3968), .VDD(VDD), .VSS(VSS), .Y(n3819) );
AND2X1 X1402 (.A(n3828), .B(n3978), .VDD(VDD), .VSS(VSS), .Y(n3829) );
AND2X1 X1403 (.A(n3838), .B(n3988), .VDD(VDD), .VSS(VSS), .Y(n3839) );
AND2X1 X1404 (.A(n3848), .B(n3998), .VDD(VDD), .VSS(VSS), .Y(n3849) );
AND2X1 X1405 (.A(N358), .B(N137), .VDD(VDD), .VSS(VSS), .Y(n3860) );
AND2X1 X1406 (.A(n3868), .B(n4018), .VDD(VDD), .VSS(VSS), .Y(n3869) );
AND2X1 X1407 (.A(n3903), .B(n4023), .VDD(VDD), .VSS(VSS), .Y(n4019) );
NOR2X1 X1408 (.A(n3725), .B(n3257), .Y(n3727), .VDD(VDD), .GND(VSS) );
NOR2X1 X1409 (.A(n3728), .B(n3561), .Y(n3725), .VDD(VDD), .GND(VSS) );
NOR2X1 X1410 (.A(n3729), .B(n3730), .Y(n3561), .VDD(VDD), .GND(VSS) );
NOR2X1 X1411 (.A(n3733), .B(n3411), .Y(n3732), .VDD(VDD), .GND(VSS) );
NOR2X1 X1412 (.A(n2228), .B(n2275), .Y(n3740), .VDD(VDD), .GND(VSS) );
NOR2X1 X1413 (.A(n3736), .B(n3742), .Y(n3738), .VDD(VDD), .GND(VSS) );
NOR2X1 X1414 (.A(n3743), .B(n2275), .Y(n3742), .VDD(VDD), .GND(VSS) );
NOR2X1 X1415 (.A(n3744), .B(n3745), .Y(n3743), .VDD(VDD), .GND(VSS) );
NOR2X1 X1416 (.A(N239), .B(n3746), .Y(n3744), .VDD(VDD), .GND(VSS) );
NOR2X1 X1417 (.A(n3721), .B(n3720), .Y(n3723), .VDD(VDD), .GND(VSS) );
NOR2X1 X1418 (.A(n3750), .B(n3751), .Y(n3715), .VDD(VDD), .GND(VSS) );
NOR2X1 X1419 (.A(n3752), .B(n3753), .Y(n3705), .VDD(VDD), .GND(VSS) );
NOR2X1 X1420 (.A(n3703), .B(n3702), .Y(n3753), .VDD(VDD), .GND(VSS) );
NOR2X1 X1421 (.A(n3754), .B(n3755), .Y(n3695), .VDD(VDD), .GND(VSS) );
NOR2X1 X1422 (.A(n3693), .B(n3692), .Y(n3755), .VDD(VDD), .GND(VSS) );
NOR2X1 X1423 (.A(n3756), .B(n3757), .Y(n3685), .VDD(VDD), .GND(VSS) );
NOR2X1 X1424 (.A(n3683), .B(n3682), .Y(n3757), .VDD(VDD), .GND(VSS) );
NOR2X1 X1425 (.A(n3758), .B(n3759), .Y(n3675), .VDD(VDD), .GND(VSS) );
NOR2X1 X1426 (.A(n3673), .B(n3672), .Y(n3759), .VDD(VDD), .GND(VSS) );
NOR2X1 X1427 (.A(n3760), .B(n3761), .Y(n3665), .VDD(VDD), .GND(VSS) );
NOR2X1 X1428 (.A(n3663), .B(n3662), .Y(n3761), .VDD(VDD), .GND(VSS) );
NOR2X1 X1429 (.A(n3762), .B(n3763), .Y(n3655), .VDD(VDD), .GND(VSS) );
NOR2X1 X1430 (.A(n3653), .B(n3652), .Y(n3763), .VDD(VDD), .GND(VSS) );
NOR2X1 X1431 (.A(n3764), .B(n3765), .Y(n3645), .VDD(VDD), .GND(VSS) );
NOR2X1 X1432 (.A(n3643), .B(n3642), .Y(n3765), .VDD(VDD), .GND(VSS) );
NOR2X1 X1433 (.A(n3766), .B(n3767), .Y(n3635), .VDD(VDD), .GND(VSS) );
NOR2X1 X1434 (.A(n3633), .B(n3632), .Y(n3767), .VDD(VDD), .GND(VSS) );
NOR2X1 X1435 (.A(n3768), .B(n3769), .Y(n3624), .VDD(VDD), .GND(VSS) );
NOR2X1 X1436 (.A(n3623), .B(n3622), .Y(n3769), .VDD(VDD), .GND(VSS) );
NOR2X1 X1437 (.A(n3772), .B(n2232), .Y(n3771), .VDD(VDD), .GND(VSS) );
NOR2X1 X1438 (.A(n3603), .B(n2271), .Y(n3623), .VDD(VDD), .GND(VSS) );
NOR2X1 X1439 (.A(n3456), .B(n2321), .Y(n3633), .VDD(VDD), .GND(VSS) );
NOR2X1 X1440 (.A(n3882), .B(n3257), .Y(n3884), .VDD(VDD), .GND(VSS) );
NOR2X1 X1441 (.A(n3885), .B(n3721), .Y(n3882), .VDD(VDD), .GND(VSS) );
NOR2X1 X1442 (.A(n3886), .B(n3887), .Y(n3721), .VDD(VDD), .GND(VSS) );
NOR2X1 X1443 (.A(n3890), .B(n3411), .Y(n3889), .VDD(VDD), .GND(VSS) );
NOR2X1 X1444 (.A(n2228), .B(n3898), .Y(n3897), .VDD(VDD), .GND(VSS) );
NOR2X1 X1445 (.A(n3878), .B(n3877), .Y(n3880), .VDD(VDD), .GND(VSS) );
NOR2X1 X1446 (.A(n3904), .B(n3905), .Y(n3872), .VDD(VDD), .GND(VSS) );
NOR2X1 X1447 (.A(n3906), .B(n3907), .Y(n3862), .VDD(VDD), .GND(VSS) );
NOR2X1 X1448 (.A(n3860), .B(n3859), .Y(n3907), .VDD(VDD), .GND(VSS) );
NOR2X1 X1449 (.A(n3908), .B(n3909), .Y(n3852), .VDD(VDD), .GND(VSS) );
NOR2X1 X1450 (.A(n3910), .B(n3911), .Y(n3842), .VDD(VDD), .GND(VSS) );
NOR2X1 X1451 (.A(n3912), .B(n3913), .Y(n3832), .VDD(VDD), .GND(VSS) );
NOR2X1 X1452 (.A(n3914), .B(n3915), .Y(n3822), .VDD(VDD), .GND(VSS) );
NOR2X1 X1453 (.A(n3916), .B(n3917), .Y(n3812), .VDD(VDD), .GND(VSS) );
NOR2X1 X1454 (.A(n3918), .B(n3919), .Y(n3802), .VDD(VDD), .GND(VSS) );
NOR2X1 X1455 (.A(n3920), .B(n3921), .Y(n3919), .VDD(VDD), .GND(VSS) );
NOR2X1 X1456 (.A(n3922), .B(n3923), .Y(n3791), .VDD(VDD), .GND(VSS) );
NOR2X1 X1457 (.A(n3924), .B(n3925), .Y(n3923), .VDD(VDD), .GND(VSS) );
NOR2X1 X1458 (.A(n3926), .B(n3927), .Y(n3781), .VDD(VDD), .GND(VSS) );
NOR2X1 X1459 (.A(n3780), .B(n3779), .Y(n3927), .VDD(VDD), .GND(VSS) );
NOR2X1 X1460 (.A(n3929), .B(n2271), .Y(n3780), .VDD(VDD), .GND(VSS) );
NAND2X1 X1461 (.A(n3578), .B(n3731), .Y(n3729), .VDD(VDD), .GND(VSS) );
NAND2X1 X1462 (.A(n3732), .B(N222), .Y(n3731), .VDD(VDD), .GND(VSS) );
NAND2X1 X1463 (.A(n3733), .B(n3734), .Y(n3578), .VDD(VDD), .GND(VSS) );
NAND2X1 X1464 (.A(N222), .B(N307), .Y(n3734), .VDD(VDD), .GND(VSS) );
NAND2X1 X1465 (.A(n3736), .B(n3737), .Y(n3735), .VDD(VDD), .GND(VSS) );
NAND2X1 X1466 (.A(n3738), .B(n3739), .Y(n3579), .VDD(VDD), .GND(VSS) );
NAND2X1 X1467 (.A(n3576), .B(N239), .Y(n3739), .VDD(VDD), .GND(VSS) );
NAND2X1 X1468 (.A(n3740), .B(n3741), .Y(n3737), .VDD(VDD), .GND(VSS) );
NAND2X1 X1469 (.A(n3612), .B(n3770), .Y(N5971), .VDD(VDD), .GND(VSS) );
NAND2X1 X1470 (.A(n3771), .B(N1), .Y(n3770), .VDD(VDD), .GND(VSS) );
NAND2X1 X1471 (.A(n3772), .B(n3773), .Y(n3612), .VDD(VDD), .GND(VSS) );
NAND2X1 X1472 (.A(N1), .B(N511), .Y(n3773), .VDD(VDD), .GND(VSS) );
NAND2X1 X1473 (.A(n3775), .B(n3776), .Y(n3613), .VDD(VDD), .GND(VSS) );
NAND2X1 X1474 (.A(n3777), .B(n3778), .Y(n3776), .VDD(VDD), .GND(VSS) );
NAND2X1 X1475 (.A(n3781), .B(n3782), .Y(n3774), .VDD(VDD), .GND(VSS) );
NAND2X1 X1476 (.A(n3787), .B(n3788), .Y(n3786), .VDD(VDD), .GND(VSS) );
NAND2X1 X1477 (.A(n3789), .B(n3790), .Y(n3787), .VDD(VDD), .GND(VSS) );
NAND2X1 X1478 (.A(n3791), .B(n3792), .Y(n3784), .VDD(VDD), .GND(VSS) );
NAND2X1 X1479 (.A(n3797), .B(n3798), .Y(n3796), .VDD(VDD), .GND(VSS) );
NAND2X1 X1480 (.A(n3799), .B(n3800), .Y(n3797), .VDD(VDD), .GND(VSS) );
NAND2X1 X1481 (.A(n3802), .B(n3803), .Y(n3794), .VDD(VDD), .GND(VSS) );
NAND2X1 X1482 (.A(n3804), .B(n3641), .Y(n3642), .VDD(VDD), .GND(VSS) );
NAND2X1 X1483 (.A(n3807), .B(n3808), .Y(n3806), .VDD(VDD), .GND(VSS) );
NAND2X1 X1484 (.A(n3809), .B(n3810), .Y(n3807), .VDD(VDD), .GND(VSS) );
NAND2X1 X1485 (.A(n3812), .B(n3813), .Y(n3804), .VDD(VDD), .GND(VSS) );
NAND2X1 X1486 (.A(n3814), .B(n3651), .Y(n3652), .VDD(VDD), .GND(VSS) );
NAND2X1 X1487 (.A(n3817), .B(n3818), .Y(n3816), .VDD(VDD), .GND(VSS) );
NAND2X1 X1488 (.A(n3819), .B(n3820), .Y(n3817), .VDD(VDD), .GND(VSS) );
NAND2X1 X1489 (.A(n3822), .B(n3823), .Y(n3814), .VDD(VDD), .GND(VSS) );
NAND2X1 X1490 (.A(n3824), .B(n3661), .Y(n3662), .VDD(VDD), .GND(VSS) );
NAND2X1 X1491 (.A(n3827), .B(n3828), .Y(n3826), .VDD(VDD), .GND(VSS) );
NAND2X1 X1492 (.A(n3829), .B(n3830), .Y(n3827), .VDD(VDD), .GND(VSS) );
NAND2X1 X1493 (.A(n3832), .B(n3833), .Y(n3824), .VDD(VDD), .GND(VSS) );
NAND2X1 X1494 (.A(n3834), .B(n3671), .Y(n3672), .VDD(VDD), .GND(VSS) );
NAND2X1 X1495 (.A(n3837), .B(n3838), .Y(n3836), .VDD(VDD), .GND(VSS) );
NAND2X1 X1496 (.A(n3839), .B(n3840), .Y(n3837), .VDD(VDD), .GND(VSS) );
NAND2X1 X1497 (.A(n3842), .B(n3843), .Y(n3834), .VDD(VDD), .GND(VSS) );
NAND2X1 X1498 (.A(n3844), .B(n3681), .Y(n3682), .VDD(VDD), .GND(VSS) );
NAND2X1 X1499 (.A(n3847), .B(n3848), .Y(n3846), .VDD(VDD), .GND(VSS) );
NAND2X1 X1500 (.A(n3849), .B(n3850), .Y(n3847), .VDD(VDD), .GND(VSS) );
NAND2X1 X1501 (.A(n3852), .B(n3853), .Y(n3844), .VDD(VDD), .GND(VSS) );
NAND2X1 X1502 (.A(n3854), .B(n3691), .Y(n3692), .VDD(VDD), .GND(VSS) );
NAND2X1 X1503 (.A(n3857), .B(n3858), .Y(n3856), .VDD(VDD), .GND(VSS) );
NAND2X1 X1504 (.A(n3862), .B(n3863), .Y(n3854), .VDD(VDD), .GND(VSS) );
NAND2X1 X1505 (.A(n3864), .B(n3701), .Y(n3702), .VDD(VDD), .GND(VSS) );
NAND2X1 X1506 (.A(n3867), .B(n3868), .Y(n3866), .VDD(VDD), .GND(VSS) );
NAND2X1 X1507 (.A(n3869), .B(n3870), .Y(n3867), .VDD(VDD), .GND(VSS) );
NAND2X1 X1508 (.A(n3872), .B(n3873), .Y(n3864), .VDD(VDD), .GND(VSS) );
NAND2X1 X1509 (.A(N171), .B(N341), .Y(n3713), .VDD(VDD), .GND(VSS) );
NAND2X1 X1510 (.A(n3880), .B(n3881), .Y(n3874), .VDD(VDD), .GND(VSS) );
NAND2X1 X1511 (.A(n3879), .B(n3749), .Y(n3881), .VDD(VDD), .GND(VSS) );
NAND2X1 X1512 (.A(N188), .B(N324), .Y(n3883), .VDD(VDD), .GND(VSS) );
NAND2X1 X1513 (.A(n3884), .B(N188), .Y(n3879), .VDD(VDD), .GND(VSS) );
NAND2X1 X1514 (.A(n3747), .B(n3888), .Y(n3886), .VDD(VDD), .GND(VSS) );
NAND2X1 X1515 (.A(n3889), .B(N205), .Y(n3888), .VDD(VDD), .GND(VSS) );
NAND2X1 X1516 (.A(n3890), .B(n3891), .Y(n3747), .VDD(VDD), .GND(VSS) );
NAND2X1 X1517 (.A(N205), .B(N307), .Y(n3891), .VDD(VDD), .GND(VSS) );
NAND2X1 X1518 (.A(n3893), .B(n3895), .Y(n3748), .VDD(VDD), .GND(VSS) );
NAND2X1 X1519 (.A(n3896), .B(n3894), .Y(n3895), .VDD(VDD), .GND(VSS) );
NAND2X1 X1520 (.A(n3899), .B(n3900), .Y(n3896), .VDD(VDD), .GND(VSS) );
NAND2X1 X1521 (.A(N273), .B(N239), .Y(n3900), .VDD(VDD), .GND(VSS) );
NAND2X1 X1522 (.A(N222), .B(N290), .Y(n3899), .VDD(VDD), .GND(VSS) );
NAND2X1 X1523 (.A(n3933), .B(n3934), .Y(n3932), .VDD(VDD), .GND(VSS) );
NAND2X1 X1524 (.A(n3937), .B(n3938), .Y(n3930), .VDD(VDD), .GND(VSS) );
NAND2X1 X1525 (.A(n3942), .B(n3943), .Y(n3941), .VDD(VDD), .GND(VSS) );
NAND2X1 X1526 (.A(n3944), .B(n3945), .Y(n3942), .VDD(VDD), .GND(VSS) );
NAND2X1 X1527 (.A(n3946), .B(n3947), .Y(n3939), .VDD(VDD), .GND(VSS) );
NAND2X1 X1528 (.A(n3951), .B(n3952), .Y(n3950), .VDD(VDD), .GND(VSS) );
NAND2X1 X1529 (.A(n3953), .B(n3954), .Y(n3951), .VDD(VDD), .GND(VSS) );
NAND2X1 X1530 (.A(n3956), .B(n3957), .Y(n3948), .VDD(VDD), .GND(VSS) );
NAND2X1 X1531 (.A(N52), .B(N443), .Y(n3810), .VDD(VDD), .GND(VSS) );
NAND2X1 X1532 (.A(n3961), .B(n3962), .Y(n3960), .VDD(VDD), .GND(VSS) );
NAND2X1 X1533 (.A(n3963), .B(n3964), .Y(n3961), .VDD(VDD), .GND(VSS) );
NAND2X1 X1534 (.A(n3966), .B(n3967), .Y(n3958), .VDD(VDD), .GND(VSS) );
NAND2X1 X1535 (.A(N69), .B(N426), .Y(n3820), .VDD(VDD), .GND(VSS) );
NAND2X1 X1536 (.A(n3971), .B(n3972), .Y(n3970), .VDD(VDD), .GND(VSS) );
NAND2X1 X1537 (.A(n3973), .B(n3974), .Y(n3971), .VDD(VDD), .GND(VSS) );
NAND2X1 X1538 (.A(n3976), .B(n3977), .Y(n3968), .VDD(VDD), .GND(VSS) );
NAND2X1 X1539 (.A(N86), .B(N409), .Y(n3830), .VDD(VDD), .GND(VSS) );
NAND2X1 X1540 (.A(n3981), .B(n3982), .Y(n3980), .VDD(VDD), .GND(VSS) );
NAND2X1 X1541 (.A(n3983), .B(n3984), .Y(n3981), .VDD(VDD), .GND(VSS) );
NAND2X1 X1542 (.A(n3986), .B(n3987), .Y(n3978), .VDD(VDD), .GND(VSS) );
NAND2X1 X1543 (.A(N103), .B(N392), .Y(n3840), .VDD(VDD), .GND(VSS) );
NAND2X1 X1544 (.A(n3991), .B(n3992), .Y(n3990), .VDD(VDD), .GND(VSS) );
NAND2X1 X1545 (.A(n3993), .B(n3994), .Y(n3991), .VDD(VDD), .GND(VSS) );
NAND2X1 X1546 (.A(n3996), .B(n3997), .Y(n3988), .VDD(VDD), .GND(VSS) );
NAND2X1 X1547 (.A(N120), .B(N375), .Y(n3850), .VDD(VDD), .GND(VSS) );
NAND2X1 X1548 (.A(n4001), .B(n4002), .Y(n4000), .VDD(VDD), .GND(VSS) );
NAND2X1 X1549 (.A(n4006), .B(n4007), .Y(n3998), .VDD(VDD), .GND(VSS) );
NAND2X1 X1550 (.A(n4008), .B(n3858), .Y(n3859), .VDD(VDD), .GND(VSS) );
NAND2X1 X1551 (.A(n4011), .B(n4012), .Y(n4010), .VDD(VDD), .GND(VSS) );
NAND2X1 X1552 (.A(n4013), .B(n4014), .Y(n4011), .VDD(VDD), .GND(VSS) );
NAND2X1 X1553 (.A(n4016), .B(n4017), .Y(n4008), .VDD(VDD), .GND(VSS) );
NAND2X1 X1554 (.A(N154), .B(N341), .Y(n3870), .VDD(VDD), .GND(VSS) );
NAND2X1 X1555 (.A(n4024), .B(n4025), .Y(n4018), .VDD(VDD), .GND(VSS) );
NAND2X1 X1556 (.A(n4023), .B(n3903), .Y(n4025), .VDD(VDD), .GND(VSS) );
NAND2X1 X1557 (.A(N171), .B(N324), .Y(n4027), .VDD(VDD), .GND(VSS) );
NAND2X1 X1558 (.A(n4028), .B(N171), .Y(n4023), .VDD(VDD), .GND(VSS) );
INVX1 X1559 (.A(N256), .AN(n2275), .VDD(VDD), .GND(VSS) );
INVX1 X1560 (.A(N511), .AN(n2232), .VDD(VDD), .GND(VSS) );
INVX1 X1561 (.A(N239), .AN(n2228), .VDD(VDD), .GND(VSS) );
INVX1 X1562 (.A(N494), .AN(n2271), .VDD(VDD), .GND(VSS) );
XOR2 X1563 (.A(n4069), .B(n3936), .Y(N5308), .VDD(VDD), .GND(VSS) );
XOR2 X1564 (.A(n3945), .B(n3944), .Y(n4071), .VDD(VDD), .GND(VSS) );
XOR2 X1565 (.A(n4066), .B(n3945), .Y(n4078), .VDD(VDD), .GND(VSS) );
XOR2 X1566 (.A(n3954), .B(n3953), .Y(n4080), .VDD(VDD), .GND(VSS) );
XOR2 X1567 (.A(n4062), .B(n3954), .Y(n4087), .VDD(VDD), .GND(VSS) );
XOR2 X1568 (.A(n3964), .B(n3963), .Y(n4089), .VDD(VDD), .GND(VSS) );
XOR2 X1569 (.A(n4095), .B(n3964), .Y(n4097), .VDD(VDD), .GND(VSS) );
XOR2 X1570 (.A(n3974), .B(n3973), .Y(n4099), .VDD(VDD), .GND(VSS) );
XOR2 X1571 (.A(n4105), .B(n3974), .Y(n4107), .VDD(VDD), .GND(VSS) );
XOR2 X1572 (.A(n3984), .B(n3983), .Y(n4109), .VDD(VDD), .GND(VSS) );
XOR2 X1573 (.A(n4115), .B(n3984), .Y(n4117), .VDD(VDD), .GND(VSS) );
XOR2 X1574 (.A(n3994), .B(n3993), .Y(n4119), .VDD(VDD), .GND(VSS) );
XOR2 X1575 (.A(n4125), .B(n3994), .Y(n4127), .VDD(VDD), .GND(VSS) );
XOR2 X1576 (.A(n4004), .B(n4003), .Y(n4129), .VDD(VDD), .GND(VSS) );
XOR2 X1577 (.A(n4003), .B(n4135), .Y(n4137), .VDD(VDD), .GND(VSS) );
XOR2 X1578 (.A(n4014), .B(n4013), .Y(n4139), .VDD(VDD), .GND(VSS) );
XOR2 X1579 (.A(n4145), .B(n4014), .Y(n4147), .VDD(VDD), .GND(VSS) );
XOR2 X1580 (.A(n4196), .B(n4076), .Y(N4946), .VDD(VDD), .GND(VSS) );
XOR2 X1581 (.A(n4085), .B(n4084), .Y(n4198), .VDD(VDD), .GND(VSS) );
XOR2 X1582 (.A(n4193), .B(n4085), .Y(n4205), .VDD(VDD), .GND(VSS) );
XOR2 X1583 (.A(n4094), .B(n4093), .Y(n4207), .VDD(VDD), .GND(VSS) );
XOR2 X1584 (.A(n4189), .B(n4094), .Y(n4214), .VDD(VDD), .GND(VSS) );
XOR2 X1585 (.A(n4104), .B(n4103), .Y(n4216), .VDD(VDD), .GND(VSS) );
XOR2 X1586 (.A(n4222), .B(n4104), .Y(n4224), .VDD(VDD), .GND(VSS) );
XOR2 X1587 (.A(n4114), .B(n4113), .Y(n4226), .VDD(VDD), .GND(VSS) );
XOR2 X1588 (.A(n4232), .B(n4114), .Y(n4234), .VDD(VDD), .GND(VSS) );
XOR2 X1589 (.A(n4124), .B(n4123), .Y(n4236), .VDD(VDD), .GND(VSS) );
XOR2 X1590 (.A(n4242), .B(n4124), .Y(n4244), .VDD(VDD), .GND(VSS) );
XOR2 X1591 (.A(n4134), .B(n4133), .Y(n4246), .VDD(VDD), .GND(VSS) );
XOR2 X1592 (.A(n4133), .B(n4252), .Y(n4254), .VDD(VDD), .GND(VSS) );
XOR2 X1593 (.A(n4144), .B(n4143), .Y(n4256), .VDD(VDD), .GND(VSS) );
XOR2 X1594 (.A(n4262), .B(n4144), .Y(n4264), .VDD(VDD), .GND(VSS) );
XOR2 X1595 (.A(n4312), .B(n4203), .Y(N4591), .VDD(VDD), .GND(VSS) );
XOR2 X1596 (.A(n4212), .B(n4211), .Y(n4314), .VDD(VDD), .GND(VSS) );
XOR2 X1597 (.A(n4309), .B(n4212), .Y(n4321), .VDD(VDD), .GND(VSS) );
OR2X1 X1598 (.A(n4075), .B(n4076), .VDD(VDD), .VSS(VSS), .Y(n4073) );
OR2X1 X1599 (.A(n4133), .B(n4134), .VDD(VDD), .VSS(VSS), .Y(n4131) );
OR2X1 X1600 (.A(n4151), .B(n4152), .VDD(VDD), .VSS(VSS), .Y(n4150) );
OR2X1 X1601 (.A(n4167), .B(n4037), .VDD(VDD), .VSS(VSS), .Y(n4166) );
OR2X1 X1602 (.A(n4202), .B(n4203), .VDD(VDD), .VSS(VSS), .Y(n4200) );
OR2X1 X1603 (.A(n4250), .B(n4251), .VDD(VDD), .VSS(VSS), .Y(n4248) );
OR2X1 X1604 (.A(n4268), .B(n4269), .VDD(VDD), .VSS(VSS), .Y(n4267) );
OR2X1 X1605 (.A(n4318), .B(n4319), .VDD(VDD), .VSS(VSS), .Y(n4316) );
AND2X1 X1606 (.A(n4031), .B(n4030), .VDD(VDD), .VSS(VSS), .Y(n4029) );
AND2X1 X1607 (.A(n3902), .B(n4036), .VDD(VDD), .VSS(VSS), .Y(n4034) );
AND2X1 X1608 (.A(n3741), .B(N222), .VDD(VDD), .VSS(VSS), .Y(n4041) );
AND2X1 X1609 (.A(n4044), .B(n4045), .VDD(VDD), .VSS(VSS), .Y(n4031) );
AND2X1 X1610 (.A(n4157), .B(n4156), .VDD(VDD), .VSS(VSS), .Y(n4021) );
AND2X1 X1611 (.A(n4014), .B(n4013), .VDD(VDD), .VSS(VSS), .Y(n4048) );
AND2X1 X1612 (.A(n4150), .B(n4149), .VDD(VDD), .VSS(VSS), .Y(n4047) );
AND2X1 X1613 (.A(n4140), .B(n4139), .VDD(VDD), .VSS(VSS), .Y(n4049) );
AND2X1 X1614 (.A(n3994), .B(n3993), .VDD(VDD), .VSS(VSS), .Y(n4052) );
AND2X1 X1615 (.A(n4130), .B(n4129), .VDD(VDD), .VSS(VSS), .Y(n4051) );
AND2X1 X1616 (.A(n3984), .B(n3983), .VDD(VDD), .VSS(VSS), .Y(n4054) );
AND2X1 X1617 (.A(n4120), .B(n4119), .VDD(VDD), .VSS(VSS), .Y(n4053) );
AND2X1 X1618 (.A(n3974), .B(n3973), .VDD(VDD), .VSS(VSS), .Y(n4056) );
AND2X1 X1619 (.A(n4110), .B(n4109), .VDD(VDD), .VSS(VSS), .Y(n4055) );
AND2X1 X1620 (.A(n3964), .B(n3963), .VDD(VDD), .VSS(VSS), .Y(n4058) );
AND2X1 X1621 (.A(n4100), .B(n4099), .VDD(VDD), .VSS(VSS), .Y(n4057) );
AND2X1 X1622 (.A(N443), .B(N35), .VDD(VDD), .VSS(VSS), .Y(n4061) );
AND2X1 X1623 (.A(n4090), .B(n4089), .VDD(VDD), .VSS(VSS), .Y(n4059) );
AND2X1 X1624 (.A(N460), .B(N18), .VDD(VDD), .VSS(VSS), .Y(n4065) );
AND2X1 X1625 (.A(n4081), .B(n4080), .VDD(VDD), .VSS(VSS), .Y(n4063) );
AND2X1 X1626 (.A(n4072), .B(n4071), .VDD(VDD), .VSS(VSS), .Y(n4067) );
AND2X1 X1627 (.A(n3934), .B(n4070), .VDD(VDD), .VSS(VSS), .Y(n4069) );
AND2X1 X1628 (.A(n3943), .B(n4079), .VDD(VDD), .VSS(VSS), .Y(n3944) );
AND2X1 X1629 (.A(n3952), .B(n4088), .VDD(VDD), .VSS(VSS), .Y(n3953) );
AND2X1 X1630 (.A(n3962), .B(n4098), .VDD(VDD), .VSS(VSS), .Y(n3963) );
AND2X1 X1631 (.A(n3972), .B(n4108), .VDD(VDD), .VSS(VSS), .Y(n3973) );
AND2X1 X1632 (.A(n3982), .B(n4118), .VDD(VDD), .VSS(VSS), .Y(n3983) );
AND2X1 X1633 (.A(n3992), .B(n4128), .VDD(VDD), .VSS(VSS), .Y(n3993) );
AND2X1 X1634 (.A(N358), .B(N120), .VDD(VDD), .VSS(VSS), .Y(n4004) );
AND2X1 X1635 (.A(n4012), .B(n4148), .VDD(VDD), .VSS(VSS), .Y(n4013) );
AND2X1 X1636 (.A(n4046), .B(n4153), .VDD(VDD), .VSS(VSS), .Y(n4149) );
AND2X1 X1637 (.A(n4161), .B(n4160), .VDD(VDD), .VSS(VSS), .Y(n4159) );
AND2X1 X1638 (.A(n4045), .B(n4166), .VDD(VDD), .VSS(VSS), .Y(n4164) );
AND2X1 X1639 (.A(N205), .B(n4170), .VDD(VDD), .VSS(VSS), .Y(n4037) );
AND2X1 X1640 (.A(n3741), .B(N188), .VDD(VDD), .VSS(VSS), .Y(n4170) );
AND2X1 X1641 (.A(n4173), .B(n4174), .VDD(VDD), .VSS(VSS), .Y(n4161) );
AND2X1 X1642 (.A(n4274), .B(n4273), .VDD(VDD), .VSS(VSS), .Y(n4151) );
AND2X1 X1643 (.A(n4144), .B(n4143), .VDD(VDD), .VSS(VSS), .Y(n4177) );
AND2X1 X1644 (.A(n4267), .B(n4266), .VDD(VDD), .VSS(VSS), .Y(n4176) );
AND2X1 X1645 (.A(n4257), .B(n4256), .VDD(VDD), .VSS(VSS), .Y(n4178) );
AND2X1 X1646 (.A(n4124), .B(n4123), .VDD(VDD), .VSS(VSS), .Y(n4181) );
AND2X1 X1647 (.A(n4247), .B(n4246), .VDD(VDD), .VSS(VSS), .Y(n4180) );
AND2X1 X1648 (.A(n4114), .B(n4113), .VDD(VDD), .VSS(VSS), .Y(n4183) );
AND2X1 X1649 (.A(n4237), .B(n4236), .VDD(VDD), .VSS(VSS), .Y(n4182) );
AND2X1 X1650 (.A(n4104), .B(n4103), .VDD(VDD), .VSS(VSS), .Y(n4185) );
AND2X1 X1651 (.A(n4227), .B(n4226), .VDD(VDD), .VSS(VSS), .Y(n4184) );
AND2X1 X1652 (.A(N426), .B(N35), .VDD(VDD), .VSS(VSS), .Y(n4188) );
AND2X1 X1653 (.A(n4217), .B(n4216), .VDD(VDD), .VSS(VSS), .Y(n4186) );
AND2X1 X1654 (.A(N443), .B(N18), .VDD(VDD), .VSS(VSS), .Y(n4192) );
AND2X1 X1655 (.A(n4208), .B(n4207), .VDD(VDD), .VSS(VSS), .Y(n4190) );
AND2X1 X1656 (.A(n4199), .B(n4198), .VDD(VDD), .VSS(VSS), .Y(n4194) );
AND2X1 X1657 (.A(n4074), .B(n4197), .VDD(VDD), .VSS(VSS), .Y(n4196) );
AND2X1 X1658 (.A(n4083), .B(n4206), .VDD(VDD), .VSS(VSS), .Y(n4084) );
AND2X1 X1659 (.A(n4092), .B(n4215), .VDD(VDD), .VSS(VSS), .Y(n4093) );
AND2X1 X1660 (.A(n4102), .B(n4225), .VDD(VDD), .VSS(VSS), .Y(n4103) );
AND2X1 X1661 (.A(n4112), .B(n4235), .VDD(VDD), .VSS(VSS), .Y(n4113) );
AND2X1 X1662 (.A(n4122), .B(n4245), .VDD(VDD), .VSS(VSS), .Y(n4123) );
AND2X1 X1663 (.A(N358), .B(N103), .VDD(VDD), .VSS(VSS), .Y(n4134) );
AND2X1 X1664 (.A(n4142), .B(n4265), .VDD(VDD), .VSS(VSS), .Y(n4143) );
AND2X1 X1665 (.A(n4175), .B(n4270), .VDD(VDD), .VSS(VSS), .Y(n4266) );
AND2X1 X1666 (.A(n4278), .B(n4277), .VDD(VDD), .VSS(VSS), .Y(n4276) );
AND2X1 X1667 (.A(n4174), .B(n4283), .VDD(VDD), .VSS(VSS), .Y(n4281) );
AND2X1 X1668 (.A(n3741), .B(N171), .VDD(VDD), .VSS(VSS), .Y(n4288) );
AND2X1 X1669 (.A(n4291), .B(n4292), .VDD(VDD), .VSS(VSS), .Y(n4278) );
AND2X1 X1670 (.A(n4261), .B(n4260), .VDD(VDD), .VSS(VSS), .Y(n4295) );
AND2X1 X1671 (.A(n4241), .B(n4240), .VDD(VDD), .VSS(VSS), .Y(n4299) );
AND2X1 X1672 (.A(n4231), .B(n4230), .VDD(VDD), .VSS(VSS), .Y(n4301) );
AND2X1 X1673 (.A(N426), .B(N18), .VDD(VDD), .VSS(VSS), .Y(n4308) );
AND2X1 X1674 (.A(n4315), .B(n4314), .VDD(VDD), .VSS(VSS), .Y(n4310) );
AND2X1 X1675 (.A(n4201), .B(n4313), .VDD(VDD), .VSS(VSS), .Y(n4312) );
NOR2X1 X1676 (.A(n4026), .B(n3257), .Y(n4028), .VDD(VDD), .GND(VSS) );
NOR2X1 X1677 (.A(n4029), .B(n3878), .Y(n4026), .VDD(VDD), .GND(VSS) );
NOR2X1 X1678 (.A(n4030), .B(n4031), .Y(n3878), .VDD(VDD), .GND(VSS) );
NOR2X1 X1679 (.A(n4034), .B(n3411), .Y(n4033), .VDD(VDD), .GND(VSS) );
NOR2X1 X1680 (.A(n4022), .B(n4021), .Y(n4024), .VDD(VDD), .GND(VSS) );
NOR2X1 X1681 (.A(n4047), .B(n4048), .Y(n4016), .VDD(VDD), .GND(VSS) );
NOR2X1 X1682 (.A(n4049), .B(n4050), .Y(n4006), .VDD(VDD), .GND(VSS) );
NOR2X1 X1683 (.A(n4004), .B(n4003), .Y(n4050), .VDD(VDD), .GND(VSS) );
NOR2X1 X1684 (.A(n4051), .B(n4052), .Y(n3996), .VDD(VDD), .GND(VSS) );
NOR2X1 X1685 (.A(n4053), .B(n4054), .Y(n3986), .VDD(VDD), .GND(VSS) );
NOR2X1 X1686 (.A(n4055), .B(n4056), .Y(n3976), .VDD(VDD), .GND(VSS) );
NOR2X1 X1687 (.A(n4057), .B(n4058), .Y(n3966), .VDD(VDD), .GND(VSS) );
NOR2X1 X1688 (.A(n4059), .B(n4060), .Y(n3956), .VDD(VDD), .GND(VSS) );
NOR2X1 X1689 (.A(n4061), .B(n4062), .Y(n4060), .VDD(VDD), .GND(VSS) );
NOR2X1 X1690 (.A(n4063), .B(n4064), .Y(n3946), .VDD(VDD), .GND(VSS) );
NOR2X1 X1691 (.A(n4065), .B(n4066), .Y(n4064), .VDD(VDD), .GND(VSS) );
NOR2X1 X1692 (.A(n4067), .B(n4068), .Y(n3937), .VDD(VDD), .GND(VSS) );
NOR2X1 X1693 (.A(n3936), .B(n3935), .Y(n4068), .VDD(VDD), .GND(VSS) );
NOR2X1 X1694 (.A(n3929), .B(n2321), .Y(n3936), .VDD(VDD), .GND(VSS) );
NOR2X1 X1695 (.A(n4156), .B(n3257), .Y(n4158), .VDD(VDD), .GND(VSS) );
NOR2X1 X1696 (.A(n4159), .B(n4022), .Y(n4156), .VDD(VDD), .GND(VSS) );
NOR2X1 X1697 (.A(n4160), .B(n4161), .Y(n4022), .VDD(VDD), .GND(VSS) );
NOR2X1 X1698 (.A(n4164), .B(n3411), .Y(n4163), .VDD(VDD), .GND(VSS) );
NOR2X1 X1699 (.A(n4152), .B(n4151), .Y(n4154), .VDD(VDD), .GND(VSS) );
NOR2X1 X1700 (.A(n4176), .B(n4177), .Y(n4146), .VDD(VDD), .GND(VSS) );
NOR2X1 X1701 (.A(n4178), .B(n4179), .Y(n4136), .VDD(VDD), .GND(VSS) );
NOR2X1 X1702 (.A(n4134), .B(n4133), .Y(n4179), .VDD(VDD), .GND(VSS) );
NOR2X1 X1703 (.A(n4180), .B(n4181), .Y(n4126), .VDD(VDD), .GND(VSS) );
NOR2X1 X1704 (.A(n4182), .B(n4183), .Y(n4116), .VDD(VDD), .GND(VSS) );
NOR2X1 X1705 (.A(n4184), .B(n4185), .Y(n4106), .VDD(VDD), .GND(VSS) );
NOR2X1 X1706 (.A(n4186), .B(n4187), .Y(n4096), .VDD(VDD), .GND(VSS) );
NOR2X1 X1707 (.A(n4188), .B(n4189), .Y(n4187), .VDD(VDD), .GND(VSS) );
NOR2X1 X1708 (.A(n4190), .B(n4191), .Y(n4086), .VDD(VDD), .GND(VSS) );
NOR2X1 X1709 (.A(n4192), .B(n4193), .Y(n4191), .VDD(VDD), .GND(VSS) );
NOR2X1 X1710 (.A(n4194), .B(n4195), .Y(n4077), .VDD(VDD), .GND(VSS) );
NOR2X1 X1711 (.A(n4076), .B(n4075), .Y(n4195), .VDD(VDD), .GND(VSS) );
NOR2X1 X1712 (.A(n3929), .B(n2377), .Y(n4076), .VDD(VDD), .GND(VSS) );
NOR2X1 X1713 (.A(n4273), .B(n3257), .Y(n4275), .VDD(VDD), .GND(VSS) );
NOR2X1 X1714 (.A(n4276), .B(n4152), .Y(n4273), .VDD(VDD), .GND(VSS) );
NOR2X1 X1715 (.A(n4277), .B(n4278), .Y(n4152), .VDD(VDD), .GND(VSS) );
NOR2X1 X1716 (.A(n4281), .B(n3411), .Y(n4280), .VDD(VDD), .GND(VSS) );
NOR2X1 X1717 (.A(n4269), .B(n4268), .Y(n4271), .VDD(VDD), .GND(VSS) );
NOR2X1 X1718 (.A(n4294), .B(n4295), .Y(n4263), .VDD(VDD), .GND(VSS) );
NOR2X1 X1719 (.A(n4296), .B(n4297), .Y(n4253), .VDD(VDD), .GND(VSS) );
NOR2X1 X1720 (.A(n4251), .B(n4250), .Y(n4297), .VDD(VDD), .GND(VSS) );
NOR2X1 X1721 (.A(n4298), .B(n4299), .Y(n4243), .VDD(VDD), .GND(VSS) );
NOR2X1 X1722 (.A(n4300), .B(n4301), .Y(n4233), .VDD(VDD), .GND(VSS) );
NOR2X1 X1723 (.A(n4302), .B(n4303), .Y(n4223), .VDD(VDD), .GND(VSS) );
NOR2X1 X1724 (.A(n4304), .B(n4305), .Y(n4303), .VDD(VDD), .GND(VSS) );
NOR2X1 X1725 (.A(n4306), .B(n4307), .Y(n4213), .VDD(VDD), .GND(VSS) );
NOR2X1 X1726 (.A(n4308), .B(n4309), .Y(n4307), .VDD(VDD), .GND(VSS) );
NOR2X1 X1727 (.A(n4310), .B(n4311), .Y(n4204), .VDD(VDD), .GND(VSS) );
NOR2X1 X1728 (.A(n4203), .B(n4202), .Y(n4311), .VDD(VDD), .GND(VSS) );
NOR2X1 X1729 (.A(n3929), .B(n2445), .Y(n4203), .VDD(VDD), .GND(VSS) );
NAND2X1 X1730 (.A(n3901), .B(n4032), .Y(n4030), .VDD(VDD), .GND(VSS) );
NAND2X1 X1731 (.A(n4033), .B(N188), .Y(n4032), .VDD(VDD), .GND(VSS) );
NAND2X1 X1732 (.A(n4034), .B(n4035), .Y(n3901), .VDD(VDD), .GND(VSS) );
NAND2X1 X1733 (.A(N188), .B(N307), .Y(n4035), .VDD(VDD), .GND(VSS) );
NAND2X1 X1734 (.A(n4037), .B(n3893), .Y(n4036), .VDD(VDD), .GND(VSS) );
NAND2X1 X1735 (.A(n4038), .B(n4039), .Y(n3902), .VDD(VDD), .GND(VSS) );
NAND2X1 X1736 (.A(n4040), .B(n3893), .Y(n4039), .VDD(VDD), .GND(VSS) );
NAND2X1 X1737 (.A(n4041), .B(N205), .Y(n3893), .VDD(VDD), .GND(VSS) );
NAND2X1 X1738 (.A(n4042), .B(n4043), .Y(n4040), .VDD(VDD), .GND(VSS) );
NAND2X1 X1739 (.A(N222), .B(N273), .Y(n4043), .VDD(VDD), .GND(VSS) );
NAND2X1 X1740 (.A(N205), .B(N290), .Y(n4042), .VDD(VDD), .GND(VSS) );
NAND2X1 X1741 (.A(n4073), .B(n4074), .Y(n4072), .VDD(VDD), .GND(VSS) );
NAND2X1 X1742 (.A(n4077), .B(n4078), .Y(n4070), .VDD(VDD), .GND(VSS) );
NAND2X1 X1743 (.A(n4082), .B(n4083), .Y(n4081), .VDD(VDD), .GND(VSS) );
NAND2X1 X1744 (.A(n4084), .B(n4085), .Y(n4082), .VDD(VDD), .GND(VSS) );
NAND2X1 X1745 (.A(n4086), .B(n4087), .Y(n4079), .VDD(VDD), .GND(VSS) );
NAND2X1 X1746 (.A(n4091), .B(n4092), .Y(n4090), .VDD(VDD), .GND(VSS) );
NAND2X1 X1747 (.A(n4093), .B(n4094), .Y(n4091), .VDD(VDD), .GND(VSS) );
NAND2X1 X1748 (.A(n4096), .B(n4097), .Y(n4088), .VDD(VDD), .GND(VSS) );
NAND2X1 X1749 (.A(N52), .B(N426), .Y(n3964), .VDD(VDD), .GND(VSS) );
NAND2X1 X1750 (.A(n4101), .B(n4102), .Y(n4100), .VDD(VDD), .GND(VSS) );
NAND2X1 X1751 (.A(n4103), .B(n4104), .Y(n4101), .VDD(VDD), .GND(VSS) );
NAND2X1 X1752 (.A(n4106), .B(n4107), .Y(n4098), .VDD(VDD), .GND(VSS) );
NAND2X1 X1753 (.A(N69), .B(N409), .Y(n3974), .VDD(VDD), .GND(VSS) );
NAND2X1 X1754 (.A(n4111), .B(n4112), .Y(n4110), .VDD(VDD), .GND(VSS) );
NAND2X1 X1755 (.A(n4113), .B(n4114), .Y(n4111), .VDD(VDD), .GND(VSS) );
NAND2X1 X1756 (.A(n4116), .B(n4117), .Y(n4108), .VDD(VDD), .GND(VSS) );
NAND2X1 X1757 (.A(N86), .B(N392), .Y(n3984), .VDD(VDD), .GND(VSS) );
NAND2X1 X1758 (.A(n4121), .B(n4122), .Y(n4120), .VDD(VDD), .GND(VSS) );
NAND2X1 X1759 (.A(n4123), .B(n4124), .Y(n4121), .VDD(VDD), .GND(VSS) );
NAND2X1 X1760 (.A(n4126), .B(n4127), .Y(n4118), .VDD(VDD), .GND(VSS) );
NAND2X1 X1761 (.A(N103), .B(N375), .Y(n3994), .VDD(VDD), .GND(VSS) );
NAND2X1 X1762 (.A(n4131), .B(n4132), .Y(n4130), .VDD(VDD), .GND(VSS) );
NAND2X1 X1763 (.A(n4136), .B(n4137), .Y(n4128), .VDD(VDD), .GND(VSS) );
NAND2X1 X1764 (.A(n4138), .B(n4002), .Y(n4003), .VDD(VDD), .GND(VSS) );
NAND2X1 X1765 (.A(n4141), .B(n4142), .Y(n4140), .VDD(VDD), .GND(VSS) );
NAND2X1 X1766 (.A(n4143), .B(n4144), .Y(n4141), .VDD(VDD), .GND(VSS) );
NAND2X1 X1767 (.A(n4146), .B(n4147), .Y(n4138), .VDD(VDD), .GND(VSS) );
NAND2X1 X1768 (.A(N137), .B(N341), .Y(n4014), .VDD(VDD), .GND(VSS) );
NAND2X1 X1769 (.A(n4154), .B(n4155), .Y(n4148), .VDD(VDD), .GND(VSS) );
NAND2X1 X1770 (.A(n4153), .B(n4046), .Y(n4155), .VDD(VDD), .GND(VSS) );
NAND2X1 X1771 (.A(N154), .B(N324), .Y(n4157), .VDD(VDD), .GND(VSS) );
NAND2X1 X1772 (.A(n4158), .B(N154), .Y(n4153), .VDD(VDD), .GND(VSS) );
NAND2X1 X1773 (.A(n4044), .B(n4162), .Y(n4160), .VDD(VDD), .GND(VSS) );
NAND2X1 X1774 (.A(n4163), .B(N171), .Y(n4162), .VDD(VDD), .GND(VSS) );
NAND2X1 X1775 (.A(n4164), .B(n4165), .Y(n4044), .VDD(VDD), .GND(VSS) );
NAND2X1 X1776 (.A(N171), .B(N307), .Y(n4165), .VDD(VDD), .GND(VSS) );
NAND2X1 X1777 (.A(n4167), .B(n4168), .Y(n4045), .VDD(VDD), .GND(VSS) );
NAND2X1 X1778 (.A(n4169), .B(n4038), .Y(n4168), .VDD(VDD), .GND(VSS) );
NAND2X1 X1779 (.A(n4171), .B(n4172), .Y(n4169), .VDD(VDD), .GND(VSS) );
NAND2X1 X1780 (.A(N205), .B(N273), .Y(n4172), .VDD(VDD), .GND(VSS) );
NAND2X1 X1781 (.A(N188), .B(N290), .Y(n4171), .VDD(VDD), .GND(VSS) );
NAND2X1 X1782 (.A(n4200), .B(n4201), .Y(n4199), .VDD(VDD), .GND(VSS) );
NAND2X1 X1783 (.A(n4204), .B(n4205), .Y(n4197), .VDD(VDD), .GND(VSS) );
NAND2X1 X1784 (.A(n4209), .B(n4210), .Y(n4208), .VDD(VDD), .GND(VSS) );
NAND2X1 X1785 (.A(n4211), .B(n4212), .Y(n4209), .VDD(VDD), .GND(VSS) );
NAND2X1 X1786 (.A(n4213), .B(n4214), .Y(n4206), .VDD(VDD), .GND(VSS) );
NAND2X1 X1787 (.A(n4218), .B(n4219), .Y(n4217), .VDD(VDD), .GND(VSS) );
NAND2X1 X1788 (.A(n4220), .B(n4221), .Y(n4218), .VDD(VDD), .GND(VSS) );
NAND2X1 X1789 (.A(n4223), .B(n4224), .Y(n4215), .VDD(VDD), .GND(VSS) );
NAND2X1 X1790 (.A(N52), .B(N409), .Y(n4104), .VDD(VDD), .GND(VSS) );
NAND2X1 X1791 (.A(n4228), .B(n4229), .Y(n4227), .VDD(VDD), .GND(VSS) );
NAND2X1 X1792 (.A(n4230), .B(n4231), .Y(n4228), .VDD(VDD), .GND(VSS) );
NAND2X1 X1793 (.A(n4233), .B(n4234), .Y(n4225), .VDD(VDD), .GND(VSS) );
NAND2X1 X1794 (.A(N69), .B(N392), .Y(n4114), .VDD(VDD), .GND(VSS) );
NAND2X1 X1795 (.A(n4238), .B(n4239), .Y(n4237), .VDD(VDD), .GND(VSS) );
NAND2X1 X1796 (.A(n4240), .B(n4241), .Y(n4238), .VDD(VDD), .GND(VSS) );
NAND2X1 X1797 (.A(n4243), .B(n4244), .Y(n4235), .VDD(VDD), .GND(VSS) );
NAND2X1 X1798 (.A(N86), .B(N375), .Y(n4124), .VDD(VDD), .GND(VSS) );
NAND2X1 X1799 (.A(n4248), .B(n4249), .Y(n4247), .VDD(VDD), .GND(VSS) );
NAND2X1 X1800 (.A(n4253), .B(n4254), .Y(n4245), .VDD(VDD), .GND(VSS) );
NAND2X1 X1801 (.A(n4255), .B(n4132), .Y(n4133), .VDD(VDD), .GND(VSS) );
NAND2X1 X1802 (.A(n4258), .B(n4259), .Y(n4257), .VDD(VDD), .GND(VSS) );
NAND2X1 X1803 (.A(n4260), .B(n4261), .Y(n4258), .VDD(VDD), .GND(VSS) );
NAND2X1 X1804 (.A(n4263), .B(n4264), .Y(n4255), .VDD(VDD), .GND(VSS) );
NAND2X1 X1805 (.A(N120), .B(N341), .Y(n4144), .VDD(VDD), .GND(VSS) );
NAND2X1 X1806 (.A(n4271), .B(n4272), .Y(n4265), .VDD(VDD), .GND(VSS) );
NAND2X1 X1807 (.A(n4270), .B(n4175), .Y(n4272), .VDD(VDD), .GND(VSS) );
NAND2X1 X1808 (.A(N137), .B(N324), .Y(n4274), .VDD(VDD), .GND(VSS) );
NAND2X1 X1809 (.A(n4275), .B(N137), .Y(n4270), .VDD(VDD), .GND(VSS) );
NAND2X1 X1810 (.A(n4173), .B(n4279), .Y(n4277), .VDD(VDD), .GND(VSS) );
NAND2X1 X1811 (.A(n4280), .B(N154), .Y(n4279), .VDD(VDD), .GND(VSS) );
NAND2X1 X1812 (.A(n4281), .B(n4282), .Y(n4173), .VDD(VDD), .GND(VSS) );
NAND2X1 X1813 (.A(N154), .B(N307), .Y(n4282), .VDD(VDD), .GND(VSS) );
NAND2X1 X1814 (.A(n4284), .B(n4167), .Y(n4283), .VDD(VDD), .GND(VSS) );
NAND2X1 X1815 (.A(n4285), .B(n4286), .Y(n4174), .VDD(VDD), .GND(VSS) );
NAND2X1 X1816 (.A(n4287), .B(n4167), .Y(n4286), .VDD(VDD), .GND(VSS) );
NAND2X1 X1817 (.A(n4288), .B(N188), .Y(n4167), .VDD(VDD), .GND(VSS) );
NAND2X1 X1818 (.A(n4289), .B(n4290), .Y(n4287), .VDD(VDD), .GND(VSS) );
NAND2X1 X1819 (.A(N188), .B(N273), .Y(n4290), .VDD(VDD), .GND(VSS) );
NAND2X1 X1820 (.A(N171), .B(N290), .Y(n4289), .VDD(VDD), .GND(VSS) );
NAND2X1 X1821 (.A(n4316), .B(n4317), .Y(n4315), .VDD(VDD), .GND(VSS) );
NAND2X1 X1822 (.A(n4320), .B(n4321), .Y(n4313), .VDD(VDD), .GND(VSS) );
INVX1 X1823 (.A(N477), .AN(n2321), .VDD(VDD), .GND(VSS) );
INVX1 X1824 (.A(N460), .AN(n2377), .VDD(VDD), .GND(VSS) );
INVX1 X1825 (.A(n4293), .AN(n4268), .VDD(VDD), .GND(VSS) );
INVX1 X1826 (.A(n4259), .AN(n4294), .VDD(VDD), .GND(VSS) );
INVX1 X1827 (.A(n4249), .AN(n4296), .VDD(VDD), .GND(VSS) );
INVX1 X1828 (.A(n4239), .AN(n4298), .VDD(VDD), .GND(VSS) );
INVX1 X1829 (.A(n4229), .AN(n4300), .VDD(VDD), .GND(VSS) );
INVX1 X1830 (.A(n4221), .AN(n4304), .VDD(VDD), .GND(VSS) );
INVX1 X1831 (.A(n4219), .AN(n4302), .VDD(VDD), .GND(VSS) );
INVX1 X1832 (.A(n4210), .AN(n4306), .VDD(VDD), .GND(VSS) );
INVX1 X1833 (.A(N443), .AN(n2445), .VDD(VDD), .GND(VSS) );
INVX1 X1834 (.A(n4309), .AN(n4211), .VDD(VDD), .GND(VSS) );
XOR2 X1835 (.A(n4221), .B(n4220), .Y(n4323), .VDD(VDD), .GND(VSS) );
XOR2 X1836 (.A(n4305), .B(n4221), .Y(n4330), .VDD(VDD), .GND(VSS) );
XOR2 X1837 (.A(n4231), .B(n4230), .Y(n4332), .VDD(VDD), .GND(VSS) );
XOR2 X1838 (.A(n4338), .B(n4231), .Y(n4340), .VDD(VDD), .GND(VSS) );
XOR2 X1839 (.A(n4241), .B(n4240), .Y(n4342), .VDD(VDD), .GND(VSS) );
XOR2 X1840 (.A(n4348), .B(n4241), .Y(n4350), .VDD(VDD), .GND(VSS) );
XOR2 X1841 (.A(n4251), .B(n4250), .Y(n4352), .VDD(VDD), .GND(VSS) );
XOR2 X1842 (.A(n4250), .B(n4358), .Y(n4360), .VDD(VDD), .GND(VSS) );
XOR2 X1843 (.A(n4261), .B(n4260), .Y(n4362), .VDD(VDD), .GND(VSS) );
XOR2 X1844 (.A(n4368), .B(n4261), .Y(n4370), .VDD(VDD), .GND(VSS) );
XOR2 X1845 (.A(n4415), .B(n4319), .Y(N4241), .VDD(VDD), .GND(VSS) );
XOR2 X1846 (.A(n4328), .B(n4327), .Y(n4417), .VDD(VDD), .GND(VSS) );
XOR2 X1847 (.A(n4412), .B(n4328), .Y(n4424), .VDD(VDD), .GND(VSS) );
XOR2 X1848 (.A(n4337), .B(n4336), .Y(n4426), .VDD(VDD), .GND(VSS) );
XOR2 X1849 (.A(n4408), .B(n4337), .Y(n4433), .VDD(VDD), .GND(VSS) );
XOR2 X1850 (.A(n4347), .B(n4346), .Y(n4435), .VDD(VDD), .GND(VSS) );
XOR2 X1851 (.A(n4441), .B(n4347), .Y(n4443), .VDD(VDD), .GND(VSS) );
XOR2 X1852 (.A(n4357), .B(n4356), .Y(n4445), .VDD(VDD), .GND(VSS) );
XOR2 X1853 (.A(n4356), .B(n4451), .Y(n4453), .VDD(VDD), .GND(VSS) );
XOR2 X1854 (.A(n4367), .B(n4366), .Y(n4455), .VDD(VDD), .GND(VSS) );
XOR2 X1855 (.A(n4461), .B(n4367), .Y(n4463), .VDD(VDD), .GND(VSS) );
XOR2 X1856 (.A(n4507), .B(n4422), .Y(N3895), .VDD(VDD), .GND(VSS) );
XOR2 X1857 (.A(n4431), .B(n4430), .Y(n4509), .VDD(VDD), .GND(VSS) );
XOR2 X1858 (.A(n4504), .B(n4431), .Y(n4516), .VDD(VDD), .GND(VSS) );
XOR2 X1859 (.A(n4440), .B(n4439), .Y(n4518), .VDD(VDD), .GND(VSS) );
XOR2 X1860 (.A(n4500), .B(n4440), .Y(n4525), .VDD(VDD), .GND(VSS) );
XOR2 X1861 (.A(n4450), .B(n4449), .Y(n4527), .VDD(VDD), .GND(VSS) );
XOR2 X1862 (.A(n4449), .B(n4533), .Y(n4535), .VDD(VDD), .GND(VSS) );
XOR2 X1863 (.A(n4460), .B(n4459), .Y(n4537), .VDD(VDD), .GND(VSS) );
XOR2 X1864 (.A(n4543), .B(n4460), .Y(n4545), .VDD(VDD), .GND(VSS) );
XOR2 X1865 (.A(n4584), .B(n4514), .Y(N3552), .VDD(VDD), .GND(VSS) );
XOR2 X1866 (.A(n4523), .B(n4522), .Y(n4586), .VDD(VDD), .GND(VSS) );
XOR2 X1867 (.A(n4581), .B(n4523), .Y(n4593), .VDD(VDD), .GND(VSS) );
XOR2 X1868 (.A(n4532), .B(n4531), .Y(n4595), .VDD(VDD), .GND(VSS) );
XOR2 X1869 (.A(n4603), .B(n4532), .Y(n4602), .VDD(VDD), .GND(VSS) );
XOR2 X1870 (.A(n4542), .B(n4541), .Y(n4605), .VDD(VDD), .GND(VSS) );
XOR2 X1871 (.A(n4611), .B(n4542), .Y(n4613), .VDD(VDD), .GND(VSS) );
OR2X1 X1872 (.A(n4356), .B(n4357), .VDD(VDD), .VSS(VSS), .Y(n4354) );
OR2X1 X1873 (.A(n4374), .B(n4375), .VDD(VDD), .VSS(VSS), .Y(n4373) );
OR2X1 X1874 (.A(n4390), .B(n4284), .VDD(VDD), .VSS(VSS), .Y(n4389) );
OR2X1 X1875 (.A(n4421), .B(n4422), .VDD(VDD), .VSS(VSS), .Y(n4419) );
OR2X1 X1876 (.A(n4449), .B(n4450), .VDD(VDD), .VSS(VSS), .Y(n4447) );
OR2X1 X1877 (.A(n4467), .B(n4468), .VDD(VDD), .VSS(VSS), .Y(n4466) );
OR2X1 X1878 (.A(n4513), .B(n4514), .VDD(VDD), .VSS(VSS), .Y(n4511) );
OR2X1 X1879 (.A(n4531), .B(n4532), .VDD(VDD), .VSS(VSS), .Y(n4529) );
OR2X1 X1880 (.A(n4549), .B(n4550), .VDD(VDD), .VSS(VSS), .Y(n4548) );
OR2X1 X1881 (.A(n4565), .B(n4483), .VDD(VDD), .VSS(VSS), .Y(n4564) );
OR2X1 X1882 (.A(n4590), .B(n4591), .VDD(VDD), .VSS(VSS), .Y(n4588) );
OR2X1 X1883 (.A(n4599), .B(n4600), .VDD(VDD), .VSS(VSS), .Y(n4597) );
AND2X1 X1884 (.A(n4219), .B(n4331), .VDD(VDD), .VSS(VSS), .Y(n4220) );
AND2X1 X1885 (.A(n4229), .B(n4341), .VDD(VDD), .VSS(VSS), .Y(n4230) );
AND2X1 X1886 (.A(n4239), .B(n4351), .VDD(VDD), .VSS(VSS), .Y(n4240) );
AND2X1 X1887 (.A(N358), .B(N86), .VDD(VDD), .VSS(VSS), .Y(n4251) );
AND2X1 X1888 (.A(n4259), .B(n4371), .VDD(VDD), .VSS(VSS), .Y(n4260) );
AND2X1 X1889 (.A(n4293), .B(n4376), .VDD(VDD), .VSS(VSS), .Y(n4372) );
AND2X1 X1890 (.A(n4384), .B(n4383), .VDD(VDD), .VSS(VSS), .Y(n4382) );
AND2X1 X1891 (.A(n4292), .B(n4389), .VDD(VDD), .VSS(VSS), .Y(n4387) );
AND2X1 X1892 (.A(N171), .B(n4393), .VDD(VDD), .VSS(VSS), .Y(n4284) );
AND2X1 X1893 (.A(n3741), .B(N154), .VDD(VDD), .VSS(VSS), .Y(n4393) );
AND2X1 X1894 (.A(n4396), .B(n4397), .VDD(VDD), .VSS(VSS), .Y(n4384) );
AND2X1 X1895 (.A(n4473), .B(n4472), .VDD(VDD), .VSS(VSS), .Y(n4374) );
AND2X1 X1896 (.A(n4367), .B(n4366), .VDD(VDD), .VSS(VSS), .Y(n4400) );
AND2X1 X1897 (.A(n4466), .B(n4465), .VDD(VDD), .VSS(VSS), .Y(n4399) );
AND2X1 X1898 (.A(n4456), .B(n4455), .VDD(VDD), .VSS(VSS), .Y(n4401) );
AND2X1 X1899 (.A(n4347), .B(n4346), .VDD(VDD), .VSS(VSS), .Y(n4404) );
AND2X1 X1900 (.A(n4446), .B(n4445), .VDD(VDD), .VSS(VSS), .Y(n4403) );
AND2X1 X1901 (.A(N392), .B(N35), .VDD(VDD), .VSS(VSS), .Y(n4407) );
AND2X1 X1902 (.A(n4436), .B(n4435), .VDD(VDD), .VSS(VSS), .Y(n4405) );
AND2X1 X1903 (.A(N409), .B(N18), .VDD(VDD), .VSS(VSS), .Y(n4411) );
AND2X1 X1904 (.A(n4427), .B(n4426), .VDD(VDD), .VSS(VSS), .Y(n4409) );
AND2X1 X1905 (.A(n4418), .B(n4417), .VDD(VDD), .VSS(VSS), .Y(n4413) );
AND2X1 X1906 (.A(n4317), .B(n4416), .VDD(VDD), .VSS(VSS), .Y(n4415) );
AND2X1 X1907 (.A(n4326), .B(n4425), .VDD(VDD), .VSS(VSS), .Y(n4327) );
AND2X1 X1908 (.A(n4335), .B(n4434), .VDD(VDD), .VSS(VSS), .Y(n4336) );
AND2X1 X1909 (.A(n4345), .B(n4444), .VDD(VDD), .VSS(VSS), .Y(n4346) );
AND2X1 X1910 (.A(N358), .B(N69), .VDD(VDD), .VSS(VSS), .Y(n4357) );
AND2X1 X1911 (.A(n4365), .B(n4464), .VDD(VDD), .VSS(VSS), .Y(n4366) );
AND2X1 X1912 (.A(n4398), .B(n4469), .VDD(VDD), .VSS(VSS), .Y(n4465) );
AND2X1 X1913 (.A(n4477), .B(n4476), .VDD(VDD), .VSS(VSS), .Y(n4475) );
AND2X1 X1914 (.A(n4397), .B(n4482), .VDD(VDD), .VSS(VSS), .Y(n4480) );
AND2X1 X1915 (.A(n3741), .B(N137), .VDD(VDD), .VSS(VSS), .Y(n4487) );
AND2X1 X1916 (.A(n4490), .B(n4491), .VDD(VDD), .VSS(VSS), .Y(n4477) );
AND2X1 X1917 (.A(n4555), .B(n4554), .VDD(VDD), .VSS(VSS), .Y(n4467) );
AND2X1 X1918 (.A(n4460), .B(n4459), .VDD(VDD), .VSS(VSS), .Y(n4494) );
AND2X1 X1919 (.A(n4548), .B(n4547), .VDD(VDD), .VSS(VSS), .Y(n4493) );
AND2X1 X1920 (.A(n4538), .B(n4537), .VDD(VDD), .VSS(VSS), .Y(n4495) );
AND2X1 X1921 (.A(N375), .B(N35), .VDD(VDD), .VSS(VSS), .Y(n4499) );
AND2X1 X1922 (.A(n4528), .B(n4527), .VDD(VDD), .VSS(VSS), .Y(n4497) );
AND2X1 X1923 (.A(N392), .B(N18), .VDD(VDD), .VSS(VSS), .Y(n4503) );
AND2X1 X1924 (.A(n4519), .B(n4518), .VDD(VDD), .VSS(VSS), .Y(n4501) );
AND2X1 X1925 (.A(n4510), .B(n4509), .VDD(VDD), .VSS(VSS), .Y(n4505) );
AND2X1 X1926 (.A(n4420), .B(n4508), .VDD(VDD), .VSS(VSS), .Y(n4507) );
AND2X1 X1927 (.A(n4429), .B(n4517), .VDD(VDD), .VSS(VSS), .Y(n4430) );
AND2X1 X1928 (.A(n4438), .B(n4526), .VDD(VDD), .VSS(VSS), .Y(n4439) );
AND2X1 X1929 (.A(N358), .B(N52), .VDD(VDD), .VSS(VSS), .Y(n4450) );
AND2X1 X1930 (.A(n4458), .B(n4546), .VDD(VDD), .VSS(VSS), .Y(n4459) );
AND2X1 X1931 (.A(n4492), .B(n4551), .VDD(VDD), .VSS(VSS), .Y(n4547) );
AND2X1 X1932 (.A(n4559), .B(n4558), .VDD(VDD), .VSS(VSS), .Y(n4557) );
AND2X1 X1933 (.A(n4491), .B(n4564), .VDD(VDD), .VSS(VSS), .Y(n4562) );
AND2X1 X1934 (.A(N137), .B(n4568), .VDD(VDD), .VSS(VSS), .Y(n4483) );
AND2X1 X1935 (.A(n3741), .B(N120), .VDD(VDD), .VSS(VSS), .Y(n4568) );
AND2X1 X1936 (.A(n4571), .B(n4572), .VDD(VDD), .VSS(VSS), .Y(n4559) );
AND2X1 X1937 (.A(n4542), .B(n4541), .VDD(VDD), .VSS(VSS), .Y(n4575) );
AND2X1 X1938 (.A(n4616), .B(n4615), .VDD(VDD), .VSS(VSS), .Y(n4574) );
AND2X1 X1939 (.A(n4606), .B(n4605), .VDD(VDD), .VSS(VSS), .Y(n4576) );
AND2X1 X1940 (.A(N375), .B(N18), .VDD(VDD), .VSS(VSS), .Y(n4580) );
AND2X1 X1941 (.A(n4596), .B(n4595), .VDD(VDD), .VSS(VSS), .Y(n4578) );
AND2X1 X1942 (.A(n4587), .B(n4586), .VDD(VDD), .VSS(VSS), .Y(n4582) );
AND2X1 X1943 (.A(n4512), .B(n4585), .VDD(VDD), .VSS(VSS), .Y(n4584) );
AND2X1 X1944 (.A(n4521), .B(n4594), .VDD(VDD), .VSS(VSS), .Y(n4522) );
AND2X1 X1945 (.A(n4530), .B(n4604), .VDD(VDD), .VSS(VSS), .Y(n4603) );
AND2X1 X1946 (.A(n4540), .B(n4614), .VDD(VDD), .VSS(VSS), .Y(n4541) );
NOR2X1 X1947 (.A(n4379), .B(n3257), .Y(n4381), .VDD(VDD), .GND(VSS) );
NOR2X1 X1948 (.A(n4382), .B(n4269), .Y(n4379), .VDD(VDD), .GND(VSS) );
NOR2X1 X1949 (.A(n4383), .B(n4384), .Y(n4269), .VDD(VDD), .GND(VSS) );
NOR2X1 X1950 (.A(n4387), .B(n3411), .Y(n4386), .VDD(VDD), .GND(VSS) );
NOR2X1 X1951 (.A(n4375), .B(n4374), .Y(n4377), .VDD(VDD), .GND(VSS) );
NOR2X1 X1952 (.A(n4399), .B(n4400), .Y(n4369), .VDD(VDD), .GND(VSS) );
NOR2X1 X1953 (.A(n4401), .B(n4402), .Y(n4359), .VDD(VDD), .GND(VSS) );
NOR2X1 X1954 (.A(n4357), .B(n4356), .Y(n4402), .VDD(VDD), .GND(VSS) );
NOR2X1 X1955 (.A(n4403), .B(n4404), .Y(n4349), .VDD(VDD), .GND(VSS) );
NOR2X1 X1956 (.A(n4405), .B(n4406), .Y(n4339), .VDD(VDD), .GND(VSS) );
NOR2X1 X1957 (.A(n4407), .B(n4408), .Y(n4406), .VDD(VDD), .GND(VSS) );
NOR2X1 X1958 (.A(n4409), .B(n4410), .Y(n4329), .VDD(VDD), .GND(VSS) );
NOR2X1 X1959 (.A(n4411), .B(n4412), .Y(n4410), .VDD(VDD), .GND(VSS) );
NOR2X1 X1960 (.A(n4413), .B(n4414), .Y(n4320), .VDD(VDD), .GND(VSS) );
NOR2X1 X1961 (.A(n4319), .B(n4318), .Y(n4414), .VDD(VDD), .GND(VSS) );
NOR2X1 X1962 (.A(n3929), .B(n2525), .Y(n4319), .VDD(VDD), .GND(VSS) );
NOR2X1 X1963 (.A(n4472), .B(n3257), .Y(n4474), .VDD(VDD), .GND(VSS) );
NOR2X1 X1964 (.A(n4475), .B(n4375), .Y(n4472), .VDD(VDD), .GND(VSS) );
NOR2X1 X1965 (.A(n4476), .B(n4477), .Y(n4375), .VDD(VDD), .GND(VSS) );
NOR2X1 X1966 (.A(n4480), .B(n3411), .Y(n4479), .VDD(VDD), .GND(VSS) );
NOR2X1 X1967 (.A(n4468), .B(n4467), .Y(n4470), .VDD(VDD), .GND(VSS) );
NOR2X1 X1968 (.A(n4493), .B(n4494), .Y(n4462), .VDD(VDD), .GND(VSS) );
NOR2X1 X1969 (.A(n4495), .B(n4496), .Y(n4452), .VDD(VDD), .GND(VSS) );
NOR2X1 X1970 (.A(n4450), .B(n4449), .Y(n4496), .VDD(VDD), .GND(VSS) );
NOR2X1 X1971 (.A(n4497), .B(n4498), .Y(n4442), .VDD(VDD), .GND(VSS) );
NOR2X1 X1972 (.A(n4499), .B(n4500), .Y(n4498), .VDD(VDD), .GND(VSS) );
NOR2X1 X1973 (.A(n4501), .B(n4502), .Y(n4432), .VDD(VDD), .GND(VSS) );
NOR2X1 X1974 (.A(n4503), .B(n4504), .Y(n4502), .VDD(VDD), .GND(VSS) );
NOR2X1 X1975 (.A(n4505), .B(n4506), .Y(n4423), .VDD(VDD), .GND(VSS) );
NOR2X1 X1976 (.A(n4422), .B(n4421), .Y(n4506), .VDD(VDD), .GND(VSS) );
NOR2X1 X1977 (.A(n3929), .B(n2617), .Y(n4422), .VDD(VDD), .GND(VSS) );
NOR2X1 X1978 (.A(n4554), .B(n3257), .Y(n4556), .VDD(VDD), .GND(VSS) );
NOR2X1 X1979 (.A(n4557), .B(n4468), .Y(n4554), .VDD(VDD), .GND(VSS) );
NOR2X1 X1980 (.A(n4558), .B(n4559), .Y(n4468), .VDD(VDD), .GND(VSS) );
NOR2X1 X1981 (.A(n4562), .B(n3411), .Y(n4561), .VDD(VDD), .GND(VSS) );
NOR2X1 X1982 (.A(n4550), .B(n4549), .Y(n4552), .VDD(VDD), .GND(VSS) );
NOR2X1 X1983 (.A(n4574), .B(n4575), .Y(n4544), .VDD(VDD), .GND(VSS) );
NOR2X1 X1984 (.A(n4576), .B(n4577), .Y(n4534), .VDD(VDD), .GND(VSS) );
NOR2X1 X1985 (.A(n4532), .B(n4531), .Y(n4577), .VDD(VDD), .GND(VSS) );
NOR2X1 X1986 (.A(n4578), .B(n4579), .Y(n4524), .VDD(VDD), .GND(VSS) );
NOR2X1 X1987 (.A(n4580), .B(n4581), .Y(n4579), .VDD(VDD), .GND(VSS) );
NOR2X1 X1988 (.A(n4582), .B(n4583), .Y(n4515), .VDD(VDD), .GND(VSS) );
NOR2X1 X1989 (.A(n4514), .B(n4513), .Y(n4583), .VDD(VDD), .GND(VSS) );
NOR2X1 X1990 (.A(n3929), .B(n2721), .Y(n4514), .VDD(VDD), .GND(VSS) );
NOR2X1 X1991 (.A(n3456), .B(n2965), .Y(n4532), .VDD(VDD), .GND(VSS) );
NAND2X1 X1992 (.A(n4322), .B(n4210), .Y(n4309), .VDD(VDD), .GND(VSS) );
NAND2X1 X1993 (.A(n4323), .B(n4324), .Y(n4210), .VDD(VDD), .GND(VSS) );
NAND2X1 X1994 (.A(n4325), .B(n4326), .Y(n4324), .VDD(VDD), .GND(VSS) );
NAND2X1 X1995 (.A(n4327), .B(n4328), .Y(n4325), .VDD(VDD), .GND(VSS) );
NAND2X1 X1996 (.A(n4329), .B(n4330), .Y(n4322), .VDD(VDD), .GND(VSS) );
NAND2X1 X1997 (.A(N35), .B(N409), .Y(n4221), .VDD(VDD), .GND(VSS) );
NAND2X1 X1998 (.A(n4332), .B(n4333), .Y(n4219), .VDD(VDD), .GND(VSS) );
NAND2X1 X1999 (.A(n4334), .B(n4335), .Y(n4333), .VDD(VDD), .GND(VSS) );
NAND2X1 X2000 (.A(n4336), .B(n4337), .Y(n4334), .VDD(VDD), .GND(VSS) );
NAND2X1 X2001 (.A(n4339), .B(n4340), .Y(n4331), .VDD(VDD), .GND(VSS) );
NAND2X1 X2002 (.A(N52), .B(N392), .Y(n4231), .VDD(VDD), .GND(VSS) );
NAND2X1 X2003 (.A(n4342), .B(n4343), .Y(n4229), .VDD(VDD), .GND(VSS) );
NAND2X1 X2004 (.A(n4344), .B(n4345), .Y(n4343), .VDD(VDD), .GND(VSS) );
NAND2X1 X2005 (.A(n4346), .B(n4347), .Y(n4344), .VDD(VDD), .GND(VSS) );
NAND2X1 X2006 (.A(n4349), .B(n4350), .Y(n4341), .VDD(VDD), .GND(VSS) );
NAND2X1 X2007 (.A(N69), .B(N375), .Y(n4241), .VDD(VDD), .GND(VSS) );
NAND2X1 X2008 (.A(n4352), .B(n4353), .Y(n4239), .VDD(VDD), .GND(VSS) );
NAND2X1 X2009 (.A(n4354), .B(n4355), .Y(n4353), .VDD(VDD), .GND(VSS) );
NAND2X1 X2010 (.A(n4359), .B(n4360), .Y(n4351), .VDD(VDD), .GND(VSS) );
NAND2X1 X2011 (.A(n4361), .B(n4249), .Y(n4250), .VDD(VDD), .GND(VSS) );
NAND2X1 X2012 (.A(n4362), .B(n4363), .Y(n4249), .VDD(VDD), .GND(VSS) );
NAND2X1 X2013 (.A(n4364), .B(n4365), .Y(n4363), .VDD(VDD), .GND(VSS) );
NAND2X1 X2014 (.A(n4366), .B(n4367), .Y(n4364), .VDD(VDD), .GND(VSS) );
NAND2X1 X2015 (.A(n4369), .B(n4370), .Y(n4361), .VDD(VDD), .GND(VSS) );
NAND2X1 X2016 (.A(N103), .B(N341), .Y(n4261), .VDD(VDD), .GND(VSS) );
NAND2X1 X2017 (.A(n4372), .B(n4373), .Y(n4259), .VDD(VDD), .GND(VSS) );
NAND2X1 X2018 (.A(n4377), .B(n4378), .Y(n4371), .VDD(VDD), .GND(VSS) );
NAND2X1 X2019 (.A(n4376), .B(n4293), .Y(n4378), .VDD(VDD), .GND(VSS) );
NAND2X1 X2020 (.A(n4379), .B(n4380), .Y(n4293), .VDD(VDD), .GND(VSS) );
NAND2X1 X2021 (.A(N120), .B(N324), .Y(n4380), .VDD(VDD), .GND(VSS) );
NAND2X1 X2022 (.A(n4381), .B(N120), .Y(n4376), .VDD(VDD), .GND(VSS) );
NAND2X1 X2023 (.A(n4291), .B(n4385), .Y(n4383), .VDD(VDD), .GND(VSS) );
NAND2X1 X2024 (.A(n4386), .B(N137), .Y(n4385), .VDD(VDD), .GND(VSS) );
NAND2X1 X2025 (.A(n4387), .B(n4388), .Y(n4291), .VDD(VDD), .GND(VSS) );
NAND2X1 X2026 (.A(N137), .B(N307), .Y(n4388), .VDD(VDD), .GND(VSS) );
NAND2X1 X2027 (.A(n4390), .B(n4391), .Y(n4292), .VDD(VDD), .GND(VSS) );
NAND2X1 X2028 (.A(n4392), .B(n4285), .Y(n4391), .VDD(VDD), .GND(VSS) );
NAND2X1 X2029 (.A(n4394), .B(n4395), .Y(n4392), .VDD(VDD), .GND(VSS) );
NAND2X1 X2030 (.A(N171), .B(N273), .Y(n4395), .VDD(VDD), .GND(VSS) );
NAND2X1 X2031 (.A(N154), .B(N290), .Y(n4394), .VDD(VDD), .GND(VSS) );
NAND2X1 X2032 (.A(n4419), .B(n4420), .Y(n4418), .VDD(VDD), .GND(VSS) );
NAND2X1 X2033 (.A(n4423), .B(n4424), .Y(n4416), .VDD(VDD), .GND(VSS) );
NAND2X1 X2034 (.A(n4428), .B(n4429), .Y(n4427), .VDD(VDD), .GND(VSS) );
NAND2X1 X2035 (.A(n4430), .B(n4431), .Y(n4428), .VDD(VDD), .GND(VSS) );
NAND2X1 X2036 (.A(n4432), .B(n4433), .Y(n4425), .VDD(VDD), .GND(VSS) );
NAND2X1 X2037 (.A(n4437), .B(n4438), .Y(n4436), .VDD(VDD), .GND(VSS) );
NAND2X1 X2038 (.A(n4439), .B(n4440), .Y(n4437), .VDD(VDD), .GND(VSS) );
NAND2X1 X2039 (.A(n4442), .B(n4443), .Y(n4434), .VDD(VDD), .GND(VSS) );
NAND2X1 X2040 (.A(N52), .B(N375), .Y(n4347), .VDD(VDD), .GND(VSS) );
NAND2X1 X2041 (.A(n4447), .B(n4448), .Y(n4446), .VDD(VDD), .GND(VSS) );
NAND2X1 X2042 (.A(n4452), .B(n4453), .Y(n4444), .VDD(VDD), .GND(VSS) );
NAND2X1 X2043 (.A(n4454), .B(n4355), .Y(n4356), .VDD(VDD), .GND(VSS) );
NAND2X1 X2044 (.A(n4457), .B(n4458), .Y(n4456), .VDD(VDD), .GND(VSS) );
NAND2X1 X2045 (.A(n4459), .B(n4460), .Y(n4457), .VDD(VDD), .GND(VSS) );
NAND2X1 X2046 (.A(n4462), .B(n4463), .Y(n4454), .VDD(VDD), .GND(VSS) );
NAND2X1 X2047 (.A(N86), .B(N341), .Y(n4367), .VDD(VDD), .GND(VSS) );
NAND2X1 X2048 (.A(n4470), .B(n4471), .Y(n4464), .VDD(VDD), .GND(VSS) );
NAND2X1 X2049 (.A(n4469), .B(n4398), .Y(n4471), .VDD(VDD), .GND(VSS) );
NAND2X1 X2050 (.A(N103), .B(N324), .Y(n4473), .VDD(VDD), .GND(VSS) );
NAND2X1 X2051 (.A(n4474), .B(N103), .Y(n4469), .VDD(VDD), .GND(VSS) );
NAND2X1 X2052 (.A(n4396), .B(n4478), .Y(n4476), .VDD(VDD), .GND(VSS) );
NAND2X1 X2053 (.A(n4479), .B(N120), .Y(n4478), .VDD(VDD), .GND(VSS) );
NAND2X1 X2054 (.A(n4480), .B(n4481), .Y(n4396), .VDD(VDD), .GND(VSS) );
NAND2X1 X2055 (.A(N120), .B(N307), .Y(n4481), .VDD(VDD), .GND(VSS) );
NAND2X1 X2056 (.A(n4483), .B(n4390), .Y(n4482), .VDD(VDD), .GND(VSS) );
NAND2X1 X2057 (.A(n4484), .B(n4485), .Y(n4397), .VDD(VDD), .GND(VSS) );
NAND2X1 X2058 (.A(n4486), .B(n4390), .Y(n4485), .VDD(VDD), .GND(VSS) );
NAND2X1 X2059 (.A(n4487), .B(N154), .Y(n4390), .VDD(VDD), .GND(VSS) );
NAND2X1 X2060 (.A(n4488), .B(n4489), .Y(n4486), .VDD(VDD), .GND(VSS) );
NAND2X1 X2061 (.A(N154), .B(N273), .Y(n4489), .VDD(VDD), .GND(VSS) );
NAND2X1 X2062 (.A(N137), .B(N290), .Y(n4488), .VDD(VDD), .GND(VSS) );
NAND2X1 X2063 (.A(n4511), .B(n4512), .Y(n4510), .VDD(VDD), .GND(VSS) );
NAND2X1 X2064 (.A(n4515), .B(n4516), .Y(n4508), .VDD(VDD), .GND(VSS) );
NAND2X1 X2065 (.A(n4520), .B(n4521), .Y(n4519), .VDD(VDD), .GND(VSS) );
NAND2X1 X2066 (.A(n4522), .B(n4523), .Y(n4520), .VDD(VDD), .GND(VSS) );
NAND2X1 X2067 (.A(n4524), .B(n4525), .Y(n4517), .VDD(VDD), .GND(VSS) );
NAND2X1 X2068 (.A(n4529), .B(n4530), .Y(n4528), .VDD(VDD), .GND(VSS) );
NAND2X1 X2069 (.A(n4534), .B(n4535), .Y(n4526), .VDD(VDD), .GND(VSS) );
NAND2X1 X2070 (.A(n4536), .B(n4448), .Y(n4449), .VDD(VDD), .GND(VSS) );
NAND2X1 X2071 (.A(n4539), .B(n4540), .Y(n4538), .VDD(VDD), .GND(VSS) );
NAND2X1 X2072 (.A(n4541), .B(n4542), .Y(n4539), .VDD(VDD), .GND(VSS) );
NAND2X1 X2073 (.A(n4544), .B(n4545), .Y(n4536), .VDD(VDD), .GND(VSS) );
NAND2X1 X2074 (.A(N69), .B(N341), .Y(n4460), .VDD(VDD), .GND(VSS) );
NAND2X1 X2075 (.A(n4552), .B(n4553), .Y(n4546), .VDD(VDD), .GND(VSS) );
NAND2X1 X2076 (.A(n4551), .B(n4492), .Y(n4553), .VDD(VDD), .GND(VSS) );
NAND2X1 X2077 (.A(N86), .B(N324), .Y(n4555), .VDD(VDD), .GND(VSS) );
NAND2X1 X2078 (.A(n4556), .B(N86), .Y(n4551), .VDD(VDD), .GND(VSS) );
NAND2X1 X2079 (.A(n4490), .B(n4560), .Y(n4558), .VDD(VDD), .GND(VSS) );
NAND2X1 X2080 (.A(n4561), .B(N103), .Y(n4560), .VDD(VDD), .GND(VSS) );
NAND2X1 X2081 (.A(n4562), .B(n4563), .Y(n4490), .VDD(VDD), .GND(VSS) );
NAND2X1 X2082 (.A(N103), .B(N307), .Y(n4563), .VDD(VDD), .GND(VSS) );
NAND2X1 X2083 (.A(n4565), .B(n4566), .Y(n4491), .VDD(VDD), .GND(VSS) );
NAND2X1 X2084 (.A(n4567), .B(n4484), .Y(n4566), .VDD(VDD), .GND(VSS) );
NAND2X1 X2085 (.A(n4569), .B(n4570), .Y(n4567), .VDD(VDD), .GND(VSS) );
NAND2X1 X2086 (.A(N137), .B(N273), .Y(n4570), .VDD(VDD), .GND(VSS) );
NAND2X1 X2087 (.A(N120), .B(N290), .Y(n4569), .VDD(VDD), .GND(VSS) );
NAND2X1 X2088 (.A(n4588), .B(n4589), .Y(n4587), .VDD(VDD), .GND(VSS) );
NAND2X1 X2089 (.A(n4592), .B(n4593), .Y(n4585), .VDD(VDD), .GND(VSS) );
NAND2X1 X2090 (.A(n4597), .B(n4598), .Y(n4596), .VDD(VDD), .GND(VSS) );
NAND2X1 X2091 (.A(n4601), .B(n4602), .Y(n4594), .VDD(VDD), .GND(VSS) );
NAND2X1 X2092 (.A(n4607), .B(n4608), .Y(n4606), .VDD(VDD), .GND(VSS) );
NAND2X1 X2093 (.A(n4609), .B(n4610), .Y(n4607), .VDD(VDD), .GND(VSS) );
NAND2X1 X2094 (.A(n4612), .B(n4613), .Y(n4604), .VDD(VDD), .GND(VSS) );
NAND2X1 X2095 (.A(N52), .B(N341), .Y(n4542), .VDD(VDD), .GND(VSS) );
INVX1 X2096 (.A(N426), .AN(n2525), .VDD(VDD), .GND(VSS) );
INVX1 X2097 (.A(N409), .AN(n2617), .VDD(VDD), .GND(VSS) );
INVX1 X2098 (.A(n4573), .AN(n4549), .VDD(VDD), .GND(VSS) );
INVX1 X2099 (.A(N392), .AN(n2721), .VDD(VDD), .GND(VSS) );
XOR2 X2100 (.A(n4651), .B(n4591), .Y(N3211), .VDD(VDD), .GND(VSS) );
XOR2 X2101 (.A(n4600), .B(n4599), .Y(n4653), .VDD(VDD), .GND(VSS) );
XOR2 X2102 (.A(n4661), .B(n4600), .Y(n4660), .VDD(VDD), .GND(VSS) );
XOR2 X2103 (.A(n4610), .B(n4609), .Y(n4663), .VDD(VDD), .GND(VSS) );
XOR2 X2104 (.A(n4646), .B(n4610), .Y(n4670), .VDD(VDD), .GND(VSS) );
XOR2 X2105 (.A(n4705), .B(n4658), .Y(N2877), .VDD(VDD), .GND(VSS) );
XOR2 X2106 (.A(n4668), .B(n4667), .Y(n4707), .VDD(VDD), .GND(VSS) );
XOR2 X2107 (.A(n4702), .B(n4668), .Y(n4714), .VDD(VDD), .GND(VSS) );
XOR2 X2108 (.A(n4746), .B(n4712), .Y(N2548), .VDD(VDD), .GND(VSS) );
OR2X1 X2109 (.A(n4657), .B(n4658), .VDD(VDD), .VSS(VSS), .Y(n4655) );
OR2X1 X2110 (.A(n4674), .B(n4675), .VDD(VDD), .VSS(VSS), .Y(n4673) );
OR2X1 X2111 (.A(n4690), .B(n4633), .VDD(VDD), .VSS(VSS), .Y(n4689) );
OR2X1 X2112 (.A(n4711), .B(n4712), .VDD(VDD), .VSS(VSS), .Y(n4709) );
OR2X1 X2113 (.A(n4718), .B(n4719), .VDD(VDD), .VSS(VSS), .Y(n4717) );
OR2X1 X2114 (.A(n4766), .B(n4734), .VDD(VDD), .VSS(VSS), .Y(n4765) );
OR2X1 X2115 (.A(n4780), .B(n4779), .VDD(VDD), .VSS(VSS), .Y(n4751) );
OR2X1 X2116 (.A(n3746), .B(n3745), .VDD(VDD), .VSS(VSS), .Y(n3898) );
AND2X1 X2117 (.A(n4573), .B(n4619), .VDD(VDD), .VSS(VSS), .Y(n4615) );
AND2X1 X2118 (.A(n4627), .B(n4626), .VDD(VDD), .VSS(VSS), .Y(n4625) );
AND2X1 X2119 (.A(n4572), .B(n4632), .VDD(VDD), .VSS(VSS), .Y(n4630) );
AND2X1 X2120 (.A(n3741), .B(N103), .VDD(VDD), .VSS(VSS), .Y(n4637) );
AND2X1 X2121 (.A(n4640), .B(n4641), .VDD(VDD), .VSS(VSS), .Y(n4627) );
AND2X1 X2122 (.A(n4680), .B(n4679), .VDD(VDD), .VSS(VSS), .Y(n4617) );
AND2X1 X2123 (.A(N341), .B(N35), .VDD(VDD), .VSS(VSS), .Y(n4645) );
AND2X1 X2124 (.A(n4673), .B(n4672), .VDD(VDD), .VSS(VSS), .Y(n4643) );
AND2X1 X2125 (.A(n4664), .B(n4663), .VDD(VDD), .VSS(VSS), .Y(n4647) );
AND2X1 X2126 (.A(n4654), .B(n4653), .VDD(VDD), .VSS(VSS), .Y(n4649) );
AND2X1 X2127 (.A(n4589), .B(n4652), .VDD(VDD), .VSS(VSS), .Y(n4651) );
AND2X1 X2128 (.A(n4598), .B(n4662), .VDD(VDD), .VSS(VSS), .Y(n4661) );
AND2X1 X2129 (.A(n4608), .B(n4671), .VDD(VDD), .VSS(VSS), .Y(n4609) );
AND2X1 X2130 (.A(n4642), .B(n4676), .VDD(VDD), .VSS(VSS), .Y(n4672) );
AND2X1 X2131 (.A(n4684), .B(n4683), .VDD(VDD), .VSS(VSS), .Y(n4682) );
AND2X1 X2132 (.A(n4641), .B(n4689), .VDD(VDD), .VSS(VSS), .Y(n4687) );
AND2X1 X2133 (.A(N103), .B(n4693), .VDD(VDD), .VSS(VSS), .Y(n4633) );
AND2X1 X2134 (.A(n3741), .B(N86), .VDD(VDD), .VSS(VSS), .Y(n4693) );
AND2X1 X2135 (.A(n4696), .B(n4697), .VDD(VDD), .VSS(VSS), .Y(n4684) );
AND2X1 X2136 (.A(n4724), .B(n4723), .VDD(VDD), .VSS(VSS), .Y(n4674) );
AND2X1 X2137 (.A(N341), .B(N18), .VDD(VDD), .VSS(VSS), .Y(n4701) );
AND2X1 X2138 (.A(n4717), .B(n4716), .VDD(VDD), .VSS(VSS), .Y(n4699) );
AND2X1 X2139 (.A(n4708), .B(n4707), .VDD(VDD), .VSS(VSS), .Y(n4703) );
AND2X1 X2140 (.A(n4656), .B(n4706), .VDD(VDD), .VSS(VSS), .Y(n4705) );
AND2X1 X2141 (.A(n4666), .B(n4715), .VDD(VDD), .VSS(VSS), .Y(n4667) );
AND2X1 X2142 (.A(n4698), .B(n4720), .VDD(VDD), .VSS(VSS), .Y(n4716) );
AND2X1 X2143 (.A(n4728), .B(n4727), .VDD(VDD), .VSS(VSS), .Y(n4726) );
AND2X1 X2144 (.A(n4697), .B(n4733), .VDD(VDD), .VSS(VSS), .Y(n4731) );
AND2X1 X2145 (.A(n3741), .B(N69), .VDD(VDD), .VSS(VSS), .Y(n4738) );
AND2X1 X2146 (.A(n4741), .B(n4742), .VDD(VDD), .VSS(VSS), .Y(n4728) );
AND2X1 X2147 (.A(n4756), .B(n4755), .VDD(VDD), .VSS(VSS), .Y(n4718) );
AND2X1 X2148 (.A(n4749), .B(n4748), .VDD(VDD), .VSS(VSS), .Y(n4744) );
AND2X1 X2149 (.A(n4710), .B(n4747), .VDD(VDD), .VSS(VSS), .Y(n4746) );
AND2X1 X2150 (.A(n4743), .B(n4752), .VDD(VDD), .VSS(VSS), .Y(n4748) );
AND2X1 X2151 (.A(n4760), .B(n4759), .VDD(VDD), .VSS(VSS), .Y(n4758) );
AND2X1 X2152 (.A(n4742), .B(n4765), .VDD(VDD), .VSS(VSS), .Y(n4763) );
AND2X1 X2153 (.A(N69), .B(n4769), .VDD(VDD), .VSS(VSS), .Y(n4734) );
AND2X1 X2154 (.A(n3741), .B(N52), .VDD(VDD), .VSS(VSS), .Y(n4769) );
AND2X1 X2155 (.A(n4772), .B(n4773), .VDD(VDD), .VSS(VSS), .Y(n4760) );
AND2X1 X2156 (.A(n4751), .B(n4750), .VDD(VDD), .VSS(VSS), .Y(n4753) );
AND2X1 X2157 (.A(n4751), .B(n4778), .VDD(VDD), .VSS(VSS), .Y(n4776) );
AND2X1 X2158 (.A(n4781), .B(n4782), .VDD(VDD), .VSS(VSS), .Y(n4779) );
AND2X1 X2159 (.A(n4773), .B(n4787), .VDD(VDD), .VSS(VSS), .Y(n4785) );
AND2X1 X2160 (.A(N18), .B(n4792), .VDD(VDD), .VSS(VSS), .Y(n4788) );
AND2X1 X2161 (.A(n4781), .B(n4799), .VDD(VDD), .VSS(VSS), .Y(n4797) );
AND2X1 X2162 (.A(N290), .B(N1), .VDD(VDD), .VSS(VSS), .Y(n4808) );
AND2X1 X2163 (.A(N545), .B(n4809), .VDD(VDD), .VSS(VSS), .Y(n4800) );
NOR2X1 X2164 (.A(n4622), .B(n3257), .Y(n4624), .VDD(VDD), .GND(VSS) );
NOR2X1 X2165 (.A(n4625), .B(n4550), .Y(n4622), .VDD(VDD), .GND(VSS) );
NOR2X1 X2166 (.A(n4626), .B(n4627), .Y(n4550), .VDD(VDD), .GND(VSS) );
NOR2X1 X2167 (.A(n4630), .B(n3411), .Y(n4629), .VDD(VDD), .GND(VSS) );
NOR2X1 X2168 (.A(n4618), .B(n4617), .Y(n4620), .VDD(VDD), .GND(VSS) );
NOR2X1 X2169 (.A(n4643), .B(n4644), .Y(n4612), .VDD(VDD), .GND(VSS) );
NOR2X1 X2170 (.A(n4645), .B(n4646), .Y(n4644), .VDD(VDD), .GND(VSS) );
NOR2X1 X2171 (.A(n4647), .B(n4648), .Y(n4601), .VDD(VDD), .GND(VSS) );
NOR2X1 X2172 (.A(n4600), .B(n4599), .Y(n4648), .VDD(VDD), .GND(VSS) );
NOR2X1 X2173 (.A(n4649), .B(n4650), .Y(n4592), .VDD(VDD), .GND(VSS) );
NOR2X1 X2174 (.A(n4591), .B(n4590), .Y(n4650), .VDD(VDD), .GND(VSS) );
NOR2X1 X2175 (.A(n3929), .B(n2837), .Y(n4591), .VDD(VDD), .GND(VSS) );
NOR2X1 X2176 (.A(n3603), .B(n2965), .Y(n4600), .VDD(VDD), .GND(VSS) );
NOR2X1 X2177 (.A(n4679), .B(n3257), .Y(n4681), .VDD(VDD), .GND(VSS) );
NOR2X1 X2178 (.A(n4682), .B(n4618), .Y(n4679), .VDD(VDD), .GND(VSS) );
NOR2X1 X2179 (.A(n4683), .B(n4684), .Y(n4618), .VDD(VDD), .GND(VSS) );
NOR2X1 X2180 (.A(n4687), .B(n3411), .Y(n4686), .VDD(VDD), .GND(VSS) );
NOR2X1 X2181 (.A(n4675), .B(n4674), .Y(n4677), .VDD(VDD), .GND(VSS) );
NOR2X1 X2182 (.A(n4699), .B(n4700), .Y(n4669), .VDD(VDD), .GND(VSS) );
NOR2X1 X2183 (.A(n4701), .B(n4702), .Y(n4700), .VDD(VDD), .GND(VSS) );
NOR2X1 X2184 (.A(n4703), .B(n4704), .Y(n4659), .VDD(VDD), .GND(VSS) );
NOR2X1 X2185 (.A(n4658), .B(n4657), .Y(n4704), .VDD(VDD), .GND(VSS) );
NOR2X1 X2186 (.A(n3929), .B(n2965), .Y(n4658), .VDD(VDD), .GND(VSS) );
NOR2X1 X2187 (.A(n4723), .B(n3257), .Y(n4725), .VDD(VDD), .GND(VSS) );
NOR2X1 X2188 (.A(n4726), .B(n4675), .Y(n4723), .VDD(VDD), .GND(VSS) );
NOR2X1 X2189 (.A(n4727), .B(n4728), .Y(n4675), .VDD(VDD), .GND(VSS) );
NOR2X1 X2190 (.A(n4731), .B(n3411), .Y(n4730), .VDD(VDD), .GND(VSS) );
NOR2X1 X2191 (.A(n4719), .B(n4718), .Y(n4721), .VDD(VDD), .GND(VSS) );
NOR2X1 X2192 (.A(n4744), .B(n4745), .Y(n4713), .VDD(VDD), .GND(VSS) );
NOR2X1 X2193 (.A(n4712), .B(n4711), .Y(n4745), .VDD(VDD), .GND(VSS) );
NOR2X1 X2194 (.A(n3929), .B(n3105), .Y(n4712), .VDD(VDD), .GND(VSS) );
NOR2X1 X2195 (.A(n4755), .B(n3257), .Y(n4757), .VDD(VDD), .GND(VSS) );
NOR2X1 X2196 (.A(n4758), .B(n4719), .Y(n4755), .VDD(VDD), .GND(VSS) );
NOR2X1 X2197 (.A(n4759), .B(n4760), .Y(n4719), .VDD(VDD), .GND(VSS) );
NOR2X1 X2198 (.A(n4763), .B(n3411), .Y(n4762), .VDD(VDD), .GND(VSS) );
NOR2X1 X2199 (.A(n4776), .B(n3257), .Y(n4775), .VDD(VDD), .GND(VSS) );
NOR2X1 X2200 (.A(n4785), .B(n3411), .Y(n4784), .VDD(VDD), .GND(VSS) );
NOR2X1 X2201 (.A(n4797), .B(n3411), .Y(n4796), .VDD(VDD), .GND(VSS) );
NOR2X1 X2202 (.A(n3898), .B(n3456), .Y(n4792), .VDD(VDD), .GND(VSS) );
NOR2X1 X2203 (.A(n4800), .B(n4806), .Y(N1581), .VDD(VDD), .GND(VSS) );
NOR2X1 X2204 (.A(n4807), .B(n4808), .Y(n4806), .VDD(VDD), .GND(VSS) );
NOR2X1 X2205 (.A(n3746), .B(n3603), .Y(n4807), .VDD(VDD), .GND(VSS) );
NOR2X1 X2206 (.A(n3929), .B(n3746), .Y(N545), .VDD(VDD), .GND(VSS) );
NOR2X1 X2207 (.A(n3745), .B(n3603), .Y(n4809), .VDD(VDD), .GND(VSS) );
NOR2X1 X2208 (.A(n3746), .B(N290), .Y(n3745), .VDD(VDD), .GND(VSS) );
NAND2X1 X2209 (.A(n4620), .B(n4621), .Y(n4614), .VDD(VDD), .GND(VSS) );
NAND2X1 X2210 (.A(n4619), .B(n4573), .Y(n4621), .VDD(VDD), .GND(VSS) );
NAND2X1 X2211 (.A(n4622), .B(n4623), .Y(n4573), .VDD(VDD), .GND(VSS) );
NAND2X1 X2212 (.A(N69), .B(N324), .Y(n4623), .VDD(VDD), .GND(VSS) );
NAND2X1 X2213 (.A(n4624), .B(N69), .Y(n4619), .VDD(VDD), .GND(VSS) );
NAND2X1 X2214 (.A(n4571), .B(n4628), .Y(n4626), .VDD(VDD), .GND(VSS) );
NAND2X1 X2215 (.A(n4629), .B(N86), .Y(n4628), .VDD(VDD), .GND(VSS) );
NAND2X1 X2216 (.A(n4630), .B(n4631), .Y(n4571), .VDD(VDD), .GND(VSS) );
NAND2X1 X2217 (.A(N86), .B(N307), .Y(n4631), .VDD(VDD), .GND(VSS) );
NAND2X1 X2218 (.A(n4633), .B(n4565), .Y(n4632), .VDD(VDD), .GND(VSS) );
NAND2X1 X2219 (.A(n4634), .B(n4635), .Y(n4572), .VDD(VDD), .GND(VSS) );
NAND2X1 X2220 (.A(n4636), .B(n4565), .Y(n4635), .VDD(VDD), .GND(VSS) );
NAND2X1 X2221 (.A(n4637), .B(N120), .Y(n4565), .VDD(VDD), .GND(VSS) );
NAND2X1 X2222 (.A(n4638), .B(n4639), .Y(n4636), .VDD(VDD), .GND(VSS) );
NAND2X1 X2223 (.A(N120), .B(N273), .Y(n4639), .VDD(VDD), .GND(VSS) );
NAND2X1 X2224 (.A(N103), .B(N290), .Y(n4638), .VDD(VDD), .GND(VSS) );
NAND2X1 X2225 (.A(n4655), .B(n4656), .Y(n4654), .VDD(VDD), .GND(VSS) );
NAND2X1 X2226 (.A(n4659), .B(n4660), .Y(n4652), .VDD(VDD), .GND(VSS) );
NAND2X1 X2227 (.A(n4665), .B(n4666), .Y(n4664), .VDD(VDD), .GND(VSS) );
NAND2X1 X2228 (.A(n4667), .B(n4668), .Y(n4665), .VDD(VDD), .GND(VSS) );
NAND2X1 X2229 (.A(n4669), .B(n4670), .Y(n4662), .VDD(VDD), .GND(VSS) );
NAND2X1 X2230 (.A(n4677), .B(n4678), .Y(n4671), .VDD(VDD), .GND(VSS) );
NAND2X1 X2231 (.A(n4676), .B(n4642), .Y(n4678), .VDD(VDD), .GND(VSS) );
NAND2X1 X2232 (.A(N52), .B(N324), .Y(n4680), .VDD(VDD), .GND(VSS) );
NAND2X1 X2233 (.A(n4681), .B(N52), .Y(n4676), .VDD(VDD), .GND(VSS) );
NAND2X1 X2234 (.A(n4640), .B(n4685), .Y(n4683), .VDD(VDD), .GND(VSS) );
NAND2X1 X2235 (.A(n4686), .B(N69), .Y(n4685), .VDD(VDD), .GND(VSS) );
NAND2X1 X2236 (.A(n4687), .B(n4688), .Y(n4640), .VDD(VDD), .GND(VSS) );
NAND2X1 X2237 (.A(N69), .B(N307), .Y(n4688), .VDD(VDD), .GND(VSS) );
NAND2X1 X2238 (.A(n4690), .B(n4691), .Y(n4641), .VDD(VDD), .GND(VSS) );
NAND2X1 X2239 (.A(n4692), .B(n4634), .Y(n4691), .VDD(VDD), .GND(VSS) );
NAND2X1 X2240 (.A(n4694), .B(n4695), .Y(n4692), .VDD(VDD), .GND(VSS) );
NAND2X1 X2241 (.A(N103), .B(N273), .Y(n4695), .VDD(VDD), .GND(VSS) );
NAND2X1 X2242 (.A(N86), .B(N290), .Y(n4694), .VDD(VDD), .GND(VSS) );
NAND2X1 X2243 (.A(n4709), .B(n4710), .Y(n4708), .VDD(VDD), .GND(VSS) );
NAND2X1 X2244 (.A(n4713), .B(n4714), .Y(n4706), .VDD(VDD), .GND(VSS) );
NAND2X1 X2245 (.A(n4721), .B(n4722), .Y(n4715), .VDD(VDD), .GND(VSS) );
NAND2X1 X2246 (.A(n4720), .B(n4698), .Y(n4722), .VDD(VDD), .GND(VSS) );
NAND2X1 X2247 (.A(N35), .B(N324), .Y(n4724), .VDD(VDD), .GND(VSS) );
NAND2X1 X2248 (.A(n4725), .B(N35), .Y(n4720), .VDD(VDD), .GND(VSS) );
NAND2X1 X2249 (.A(n4696), .B(n4729), .Y(n4727), .VDD(VDD), .GND(VSS) );
NAND2X1 X2250 (.A(n4730), .B(N52), .Y(n4729), .VDD(VDD), .GND(VSS) );
NAND2X1 X2251 (.A(n4731), .B(n4732), .Y(n4696), .VDD(VDD), .GND(VSS) );
NAND2X1 X2252 (.A(N52), .B(N307), .Y(n4732), .VDD(VDD), .GND(VSS) );
NAND2X1 X2253 (.A(n4734), .B(n4690), .Y(n4733), .VDD(VDD), .GND(VSS) );
NAND2X1 X2254 (.A(n4735), .B(n4736), .Y(n4697), .VDD(VDD), .GND(VSS) );
NAND2X1 X2255 (.A(n4737), .B(n4690), .Y(n4736), .VDD(VDD), .GND(VSS) );
NAND2X1 X2256 (.A(n4738), .B(N86), .Y(n4690), .VDD(VDD), .GND(VSS) );
NAND2X1 X2257 (.A(n4739), .B(n4740), .Y(n4737), .VDD(VDD), .GND(VSS) );
NAND2X1 X2258 (.A(N86), .B(N273), .Y(n4740), .VDD(VDD), .GND(VSS) );
NAND2X1 X2259 (.A(N69), .B(N290), .Y(n4739), .VDD(VDD), .GND(VSS) );
NAND2X1 X2260 (.A(n4750), .B(n4751), .Y(n4749), .VDD(VDD), .GND(VSS) );
NAND2X1 X2261 (.A(n4753), .B(n4754), .Y(n4747), .VDD(VDD), .GND(VSS) );
NAND2X1 X2262 (.A(n4752), .B(n4743), .Y(n4754), .VDD(VDD), .GND(VSS) );
NAND2X1 X2263 (.A(N18), .B(N324), .Y(n4756), .VDD(VDD), .GND(VSS) );
NAND2X1 X2264 (.A(n4757), .B(N18), .Y(n4752), .VDD(VDD), .GND(VSS) );
NAND2X1 X2265 (.A(n4741), .B(n4761), .Y(n4759), .VDD(VDD), .GND(VSS) );
NAND2X1 X2266 (.A(n4762), .B(N35), .Y(n4761), .VDD(VDD), .GND(VSS) );
NAND2X1 X2267 (.A(n4763), .B(n4764), .Y(n4741), .VDD(VDD), .GND(VSS) );
NAND2X1 X2268 (.A(N35), .B(N307), .Y(n4764), .VDD(VDD), .GND(VSS) );
NAND2X1 X2269 (.A(n4766), .B(n4767), .Y(n4742), .VDD(VDD), .GND(VSS) );
NAND2X1 X2270 (.A(n4768), .B(n4735), .Y(n4767), .VDD(VDD), .GND(VSS) );
NAND2X1 X2271 (.A(n4770), .B(n4771), .Y(n4768), .VDD(VDD), .GND(VSS) );
NAND2X1 X2272 (.A(N69), .B(N273), .Y(n4771), .VDD(VDD), .GND(VSS) );
NAND2X1 X2273 (.A(N52), .B(N290), .Y(n4770), .VDD(VDD), .GND(VSS) );
NAND2X1 X2274 (.A(n4750), .B(n4774), .Y(N2223), .VDD(VDD), .GND(VSS) );
NAND2X1 X2275 (.A(n4775), .B(N1), .Y(n4774), .VDD(VDD), .GND(VSS) );
NAND2X1 X2276 (.A(n4776), .B(n4777), .Y(n4750), .VDD(VDD), .GND(VSS) );
NAND2X1 X2277 (.A(N1), .B(N324), .Y(n4777), .VDD(VDD), .GND(VSS) );
NAND2X1 X2278 (.A(n4779), .B(n4780), .Y(n4778), .VDD(VDD), .GND(VSS) );
NAND2X1 X2279 (.A(n4772), .B(n4783), .Y(n4780), .VDD(VDD), .GND(VSS) );
NAND2X1 X2280 (.A(n4784), .B(N18), .Y(n4783), .VDD(VDD), .GND(VSS) );
NAND2X1 X2281 (.A(n4785), .B(n4786), .Y(n4772), .VDD(VDD), .GND(VSS) );
NAND2X1 X2282 (.A(N18), .B(N307), .Y(n4786), .VDD(VDD), .GND(VSS) );
NAND2X1 X2283 (.A(n4788), .B(n4766), .Y(n4787), .VDD(VDD), .GND(VSS) );
NAND2X1 X2284 (.A(n4789), .B(n4790), .Y(n4773), .VDD(VDD), .GND(VSS) );
NAND2X1 X2285 (.A(n4791), .B(n4766), .Y(n4790), .VDD(VDD), .GND(VSS) );
NAND2X1 X2286 (.A(n4792), .B(N52), .Y(n4766), .VDD(VDD), .GND(VSS) );
NAND2X1 X2287 (.A(n4793), .B(n4794), .Y(n4791), .VDD(VDD), .GND(VSS) );
NAND2X1 X2288 (.A(N52), .B(N273), .Y(n4794), .VDD(VDD), .GND(VSS) );
NAND2X1 X2289 (.A(N35), .B(N290), .Y(n4793), .VDD(VDD), .GND(VSS) );
NAND2X1 X2290 (.A(n4782), .B(n4795), .Y(N1901), .VDD(VDD), .GND(VSS) );
NAND2X1 X2291 (.A(n4796), .B(N1), .Y(n4795), .VDD(VDD), .GND(VSS) );
NAND2X1 X2292 (.A(n4797), .B(n4798), .Y(n4782), .VDD(VDD), .GND(VSS) );
NAND2X1 X2293 (.A(N1), .B(N307), .Y(n4798), .VDD(VDD), .GND(VSS) );
NAND2X1 X2294 (.A(n4800), .B(n4789), .Y(n4799), .VDD(VDD), .GND(VSS) );
NAND2X1 X2295 (.A(n4801), .B(n4802), .Y(n4781), .VDD(VDD), .GND(VSS) );
NAND2X1 X2296 (.A(n4803), .B(n4789), .Y(n4802), .VDD(VDD), .GND(VSS) );
NAND2X1 X2297 (.A(n4804), .B(n4805), .Y(n4803), .VDD(VDD), .GND(VSS) );
NAND2X1 X2298 (.A(N35), .B(N273), .Y(n4805), .VDD(VDD), .GND(VSS) );
NAND2X1 X2299 (.A(N18), .B(N290), .Y(n4804), .VDD(VDD), .GND(VSS) );
INVX1 X2300 (.A(N375), .AN(n2837), .VDD(VDD), .GND(VSS) );
INVX1 X2301 (.A(N358), .AN(n2965), .VDD(VDD), .GND(VSS) );
INVX1 X2302 (.A(N341), .AN(n3105), .VDD(VDD), .GND(VSS) );
INVX1 X2303 (.A(N324), .AN(n3257), .VDD(VDD), .GND(VSS) );
INVX1 X2304 (.A(N307), .AN(n3411), .VDD(VDD), .GND(VSS) );
INVX1 X2305 (.A(N35), .AN(n3456), .VDD(VDD), .GND(VSS) );
INVX1 X2306 (.A(N1), .AN(n3929), .VDD(VDD), .GND(VSS) );
INVX1 X2307 (.A(N18), .AN(n3603), .VDD(VDD), .GND(VSS) );
OR2X1 X2308 (.A(n4617), .B(n4618), .VDD(VDD), .VSS(VSS), .Y(n4616) );
AND2X1 X2309 (.A(n2505), .B(n2504), .VDD(VDD), .VSS(VSS), .Y(n2533) );
NAND2X1 X2310 (.A(n2838), .B(n2839), .Y(n2724), .VDD(VDD), .GND(VSS) );
NAND2X1 X2311 (.A(n3139), .B(n3140), .Y(n3137), .VDD(VDD), .GND(VSS) );
INVX1 X2312 (.A(N273), .AN(n3746), .VDD(VDD), .GND(VSS) );

endmodule 
//////////////////////////////////

