.SUBCKT c432 N1 N4 N8 N11 N14 N17 N21 N24 N27 N30 N34 N37 N40 N43 N47 N50 N53 N56 N60 N63 N66 N69 N73 N76 N79 N82 N86 N89 N92 N95 N99 N102 N105 N108 N112 N115 N223 N329 N370 N421 N430 N431 N432 VDD VSS 
M1 N432 n178 VDD VDD pmos w=2u l=1u
M2 N432 n179 VDD VDD pmos w=2u l=1u
M3 net n178 GND GND nmos w=1u l=1u
M4 N432 n179 net GND nmos w=1u l=1u
M5 n179 n181 n0 GND nmos w=1u l=1u
M6 n0 n180 GND GND nmos w=1u l=1u 
M7 n179 n181 VDD VDD pmos w=2u l=1u
M8 n179 n180 VDD VDD pmos w=2u l=1u
M9 n180 n183 VDD VDD pmos w=2u l=1u
M10 n180 n182 VDD VDD pmos w=2u l=1u
M11 n180 n183 n0 VSS nmos w=1u l=1u
M12 n0 n182 VSS VSS nmos w=1u l=1u 
M13 n0 n185 net VDD pmos w=2u l=1u
M14 n183 n0 VDD VDD pmos w=2u l=1u
M15 net n184 VDD VDD pmos w=2u l=1u
M16 n183 n0 VSS VSS nmos w=1u l=1u
M17 n0 n184 VSS VSS nmos w=1u l=1u
M18 n0 n185 VSS VSS nmos w=1u l=1u
M19 n182 n187 net41 VDD pmos w=2u l=1u
M20 net41 n186 VDD VDD pmos w=2u l=1u
M21 n182 n187 GND GND nmos w=1u l=1u
M22 n182 n186 GND GND nmos w=1u l=1u 
M23 n187 n189 net41 VDD pmos w=2u l=1u  
M24 net41 n188 VDD VDD pmos w=2u l=1u
M25 n187 n189 GND GND nmos w=1u l=1u
M26 n187 n188 GND GND nmos w=1u l=1u
M27 n186 n191 GND GND nmos w=1u l=1u
M28 n186 n190 GND GND nmos w=1u l=1u
M29 n186 n191 net41 VDD pmos w=2u l=1u
M30 net41 n190 VDD VDD pmos w=2u l=1u
M31 n190 n193 GND GND nmos w=1u l=1u
M32 n190 n192 GND GND nmos w=1u l=1u
M33 n190 n193 net41 VDD pmos w=2u l=1u
M34 net41 n192 VDD VDD pmos w=2u l=1u
M35 n192 n194 GND GND nmos w=1u l=1u
M36 n192 N329 GND GND nmos w=1u l=1u
M37 n192 n194 net41 VDD pmos w=2u l=1u 
M38 net41 N329 VDD VDD pmos w=2u l=1u
M39 N431 n196 n0 GND nmos w=1u l=1u
M40 n0 n195 GND GND nmos w=1u l=1u
M41 N431 n196 VDD VDD pmos w=2u l=1u
M42 N431 n195 VDD VDD pmos w=2u l=1u
M43 n196 n198 n0 GND nmos w=1u l=1u
M44 n0 n197 GND GND nmos w=1u l=1u
M45 n196 n198 VDD VDD pmos w=2u l=1u
M46 n196 n197 VDD VDD pmos w=2u l=1u 
M47 n197 n199 GND GND nmos w=1u l=1u
M48 n197 n185 GND GND nmos w=1u l=1u
M49 n197 n199 net41 VDD pmos w=2u l=1u 
M50 net41 n185 VDD VDD pmos w=2u l=1u
M51 n195 n201 GND GND nmos w=1u l=1u
M52 n195 n200 GND GND nmos w=1u l=1u
M53 n195 n201 net41 VDD pmos w=2u l=1u
M54 net41 n200 VDD VDD pmos w=2u l=1u
M55 N421 n203 GND GND nmos w=1u l=1u
M56 N421 n202 GND GND nmos w=1u l=1u
M57 N421 n203 net41 VDD pmos w=2u l=1u
M58 net41 n202 VDD VDD pmos w=2u l=1u
M59 n203 n205 GND GND nmos w=1u l=1u
M60 n203 n204 GND GND nmos w=1u l=1u
M61 n203 n205 net41 VDD pmos w=2u l=1u
M62 net41 n204 VDD VDD pmos w=2u l=1u
M63 n205 n189 n0 GND nmos w=1u l=1u
M64 n0 n206 GND GND nmos w=1u l=1u
M65 n205 n189 VDD VDD pmos w=2u l=1u
M66 n205 n206 VDD VDD pmos w=2u l=1u
M67 n189 n208 n0 GND nmos w=1u l=1u
M68 n0 n207 GND GND nmos w=1u l=1u
M69 n189 n208 VDD VDD pmos w=2u l=1u
M70 n189 n207 VDD VDD pmos w=2u l=1u
M71 n207 n210 GND GND nmos w=1u l=1u
M72 n207 n209 GND GND nmos w=1u l=1u
M73 n207 n210 net41 VDD pmos w=2u l=1u
M74 net41 n209 VDD VDD pmos w=2u l=1u
M75 n210 n212 GND GND nmos w=1u l=1u
M76 n210 n211 GND GND nmos w=1u l=1u
M77 n210 n212 net41 VDD pmos w=2u l=1u
M78 net41 n211 VDD VDD pmos w=2u l=1u
M79 n209 n214 GND GND nmos w=1u l=1u
M80 n209 n213 GND GND nmos w=1u l=1u
M81 n209 n214 net41 VDD pmos w=2u l=1u
M82 net41 n213 VDD VDD pmos w=2u l=1u
M83 n206 n198 VDD VDD pmos w=2u l=1u
M84 n206 n198 GND GND nmos w=1u l=1u
M85 n198 n215 n0 GND nmos w=1u l=1u
M86 n0 n184 GND GND nmos w=1u l=1u
M87 n198 n215 VDD VDD pmos w=2u l=1u
M88 n198 n184 VDD VDD pmos w=2u l=1u
M89 n215 n188 VDD VDD pmos w=2u l=1u
M90 n215 n188 GND GND nmos w=1u l=1u
M91 n188 n217 GND GND nmos w=1u l=1u
M92 n188 n216 GND GND nmos w=1u l=1u
M93 n188 n217 net41 VDD pmos w=2u l=1u
M94 net41 n216 VDD VDD pmos w=2u l=1u
M95 n216 n0 GND GND nmos w=1u l=1u
M96 n0 n218 GND GND nmos w=1u l=1u
M97 n0 n219 GND GND nmos w=1u l=1u
M98 n0 n219 n1 VDD pmos w=2u l=1u
M99 n216 n0 VDD VDD pmos w=2u l=1u
M100 n1 n218 VDD VDD pmos w=2u l=1u
M101 n219 n220 GND GND nmos w=1u l=1u
M102 n219 n211 GND GND nmos w=1u l=1u
M103 n219 n220 net41 VDD pmos w=2u l=1u
M104 net41 n211 VDD VDD pmos w=2u l=1u
M105 n218 n0 GND GND nmos w=1u l=1u
M106 net127 N86 GND GND nmos w=1u l=1u
M107 n0 N329 net127 GND nmos w=1u l=1u
M108 n0 N86 VDD VDD pmos w=2u l=1u
M109 n0 N329 VDD VDD pmos w=2u l=1u
M110 n218 n0 VDD VDD pmos w=2u l=1u
M111 n184 n222 n0 GND nmos w=1u l=1u
M112 n0 n221 GND GND nmos w=1u l=1u
M113 n184 n222 VDD VDD pmos w=2u l=1u
M114 n184 n221 VDD VDD pmos w=2u l=1u
M115 n221 n224 GND GND nmos w=1u l=1u
M116 n221 n223 GND GND nmos w=1u l=1u
M117 n221 n224 net41 VDD pmos w=2u l=1u
M118 net41 n223 VDD VDD pmos w=2u l=1u
M119 n224 n0 GND GND nmos w=1u l=1u
M120 net127 N79 GND GND nmos w=1u l=1u
M121 n0 N370 net127 GND nmos w=1u l=1u
M122 n0 N79 VDD VDD pmos w=2u l=1u
M123 n0 N370 VDD VDD pmos w=2u l=1u
M124 n224 n0 VDD VDD pmos w=2u l=1u
M125 n223 n225 GND GND nmos w=1u l=1u
M126 n223 n213 GND GND nmos w=1u l=1u
M127 n223 n225 net41 VDD pmos w=2u l=1u
M128 net41 n213 VDD VDD pmos w=2u l=1u
M129 n204 n0 GND GND nmos w=1u l=1u
M130 n0 N430 GND GND nmos w=1u l=1u
M131 n0 N108 GND GND nmos w=1u l=1u
M132 n0 N108 n1 VDD pmos w=2u l=1u
M133 n204 n0 VDD VDD pmos w=2u l=1u
M134 n1 N430 VDD VDD pmos w=2u l=1u
M135 N430 n227 n0 GND nmos w=1u l=1u
M136 n0 n226 GND GND nmos w=1u l=1u
M137 N430 n227 VDD VDD pmos w=2u l=1u
M138 N430 n226 VDD VDD pmos w=2u l=1u
M139 n227 n200 GND GND nmos w=1u l=1u
M140 n227 n185 GND GND nmos w=1u l=1u
M141 n227 n200 net41 VDD pmos w=2u l=1u
M142 net41 n185 VDD VDD pmos w=2u l=1u
M143 n200 n178 VDD VDD pmos w=2u l=1u
M144 n200 n178 GND GND nmos w=1u l=1u
M145 n178 n229 n0 GND nmos w=1u l=1u
M146 n0 n228 GND GND nmos w=1u l=1u
M147 n178 n229 VDD VDD pmos w=2u l=1u
M148 n178 n228 VDD VDD pmos w=2u l=1u
M149 n228 n231 GND GND nmos w=1u l=1u
M150 n228 n230 GND GND nmos w=1u l=1u
M151 n228 n231 net41 VDD pmos w=2u l=1u
M152 net41 n230 VDD VDD pmos w=2u l=1u
M153 n231 n0 GND GND nmos w=1u l=1u
M154 net127 N27 GND GND nmos w=1u l=1u
M155 n0 N370 net127 GND nmos w=1u l=1u
M156 n0 N27 VDD VDD pmos w=2u l=1u
M157 n0 N370 VDD VDD pmos w=2u l=1u
M158 n231 n0 VDD VDD pmos w=2u l=1u
M159 n230 n232 GND GND nmos w=1u l=1u
M160 n230 n213 GND GND nmos w=1u l=1u
M161 n230 n232 net41 VDD pmos w=2u l=1u
M162 net41 n213 VDD VDD pmos w=2u l=1u
M163 n185 n0 GND GND nmos w=1u l=1u
M164 net127 n234 GND GND nmos w=1u l=1u
M165 n0 n233 net127 GND nmos w=1u l=1u
M166 n0 n234 VDD VDD pmos w=2u l=1u
M167 n0 n233 VDD VDD pmos w=2u l=1u
M168 n185 n0 VDD VDD pmos w=2u l=1u
M169 n233 n236 GND GND nmos w=1u l=1u
M170 n233 n235 GND GND nmos w=1u l=1u
M171 n233 n236 net41 VDD pmos w=2u l=1u
M172 net41 n235 VDD VDD pmos w=2u l=1u
M173 n236 n237 GND GND nmos w=1u l=1u
M174 n236 n213 GND GND nmos w=1u l=1u
M175 n236 n237 net41 VDD pmos w=2u l=1u
M176 net41 n213 VDD VDD pmos w=2u l=1u
M177 n235 n0 GND GND nmos w=1u l=1u
M178 net127 N66 GND GND nmos w=1u l=1u
M179 n0 N370 net127 GND nmos w=1u l=1u
M180 n0 N66 VDD VDD pmos w=2u l=1u
M181 n0 N370 VDD VDD pmos w=2u l=1u
M182 n235 n0 VDD VDD pmos w=2u l=1u
M183 n226 n199 GND GND nmos w=1u l=1u
M184 n226 n201 GND GND nmos w=1u l=1u
M185 n226 n199 net41 VDD pmos w=2u l=1u
M186 net41 n201 VDD VDD pmos w=2u l=1u
M187 n199 n0 GND GND nmos w=1u l=1u
M188 net127 n239 GND GND nmos w=1u l=1u
M189 n0 n238 net127 GND nmos w=1u l=1u
M190 n0 n239 VDD VDD pmos w=2u l=1u
M191 n0 n238 VDD VDD pmos w=2u l=1u
M192 n199 n0 VDD VDD pmos w=2u l=1u
M193 n238 n191 GND GND nmos w=1u l=1u
M194 n238 n240 GND GND nmos w=1u l=1u
M195 n238 n191 net41 VDD pmos w=2u l=1u
M196 net41 n240 VDD VDD pmos w=2u l=1u
M197 n191 n241 GND GND nmos w=1u l=1u
M198 n191 n211 GND GND nmos w=1u l=1u
M199 n191 n241 net41 VDD pmos w=2u l=1u
M200 net41 n211 VDD VDD pmos w=2u l=1u
M201 n241 N53 VDD VDD pmos w=2u l=1u
M202 n241 N53 GND GND nmos w=1u l=1u
M203 n211 N370 VDD VDD pmos w=2u l=1u
M204 n211 N370 GND GND nmos w=1u l=1u
M205 n240 n0 GND GND nmos w=1u l=1u
M206 net127 N47 GND GND nmos w=1u l=1u
M207 n0 N329 net127 GND nmos w=1u l=1u
M208 n0 N47 VDD VDD pmos w=2u l=1u
M209 n0 N329 VDD VDD pmos w=2u l=1u
M210 n240 n0 VDD VDD pmos w=2u l=1u
M211 n201 n181 VDD VDD pmos w=2u l=1u
M212 n201 n181 GND GND nmos w=1u l=1u
M213 n181 n243 n0 GND nmos w=1u l=1u
M214 n0 n242 GND GND nmos w=1u l=1u
M215 n181 n243 VDD VDD pmos w=2u l=1u
M216 n181 n242 VDD VDD pmos w=2u l=1u
M217 n243 n245 GND GND nmos w=1u l=1u
M218 n243 n244 GND GND nmos w=1u l=1u
M219 n243 n245 net41 VDD pmos w=2u l=1u
M220 net41 n244 VDD VDD pmos w=2u l=1u
M221 n245 n0 GND GND nmos w=1u l=1u
M222 net127 N34 GND GND nmos w=1u l=1u
M223 n0 N329 net127 GND nmos w=1u l=1u
M224 n0 N34 VDD VDD pmos w=2u l=1u
M225 n0 N329 VDD VDD pmos w=2u l=1u
M226 n245 n0 VDD VDD pmos w=2u l=1u
M227 n242 n247 GND GND nmos w=1u l=1u
M228 n242 n246 GND GND nmos w=1u l=1u
M229 n242 n247 net41 VDD pmos w=2u l=1u
M230 net41 n246 VDD VDD pmos w=2u l=1u
M231 n246 n0 GND GND nmos w=1u l=1u
M232 net127 N40 GND GND nmos w=1u l=1u
M233 n0 N370 net127 GND nmos w=1u l=1u
M234 n0 N40 VDD VDD pmos w=2u l=1u
M235 n0 N370 VDD VDD pmos w=2u l=1u
M236 n246 n0 VDD VDD pmos w=2u l=1u
M237 n202 n249 GND GND nmos w=1u l=1u
M238 n202 n248 GND GND nmos w=1u l=1u
M239 n202 n249 net41 VDD pmos w=2u l=1u
M240 net41 n248 VDD VDD pmos w=2u l=1u
M241 n249 n250 n0 GND nmos w=1u l=1u
M242 n0 N4 GND GND nmos w=1u l=1u
M243 n249 n250 VDD VDD pmos w=2u l=1u
M244 n249 N4 VDD VDD pmos w=2u l=1u
M245 n250 N370 n0 GND nmos w=1u l=1u
M246 n0 N14 GND GND nmos w=1u l=1u
M247 n250 N370 VDD VDD pmos w=2u l=1u
M248 n250 N14 VDD VDD pmos w=2u l=1u
M249 n248 n252 n0 GND nmos w=1u l=1u
M250 n0 n251 GND GND nmos w=1u l=1u
M251 n248 n252 VDD VDD pmos w=2u l=1u
M252 n248 n251 VDD VDD pmos w=2u l=1u
M253 n251 N329 n0 GND nmos w=1u l=1u
M254 n0 N8 GND GND nmos w=1u l=1u
M255 n251 N329 VDD VDD pmos w=2u l=1u
M256 n251 N8 VDD VDD pmos w=2u l=1u
M257 N370 n254 n0 GND nmos w=1u l=1u
M258 n0 n253 GND GND nmos w=1u l=1u
M259 N370 n254 VDD VDD pmos w=2u l=1u
M260 N370 n253 VDD VDD pmos w=2u l=1u
M261 n254 n256 GND GND nmos w=1u l=1u
M262 n254 n255 GND GND nmos w=1u l=1u
M263 n254 n256 net41 VDD pmos w=2u l=1u
M264 net41 n255 VDD VDD pmos w=2u l=1u
M265 n256 n258 n0 GND nmos w=1u l=1u
M266 n0 n257 GND GND nmos w=1u l=1u
M267 n256 n258 VDD VDD pmos w=2u l=1u
M268 n256 n257 VDD VDD pmos w=2u l=1u
M269 n258 n260 n0 GND nmos w=1u l=1u
M270 n0 n259 GND GND nmos w=1u l=1u
M271 n258 n260 VDD VDD pmos w=2u l=1u
M272 n258 n259 VDD VDD pmos w=2u l=1u
M273 n260 n261 VDD VDD pmos w=2u l=1u
M274 n260 n261 GND GND nmos w=1u l=1u
M275 n259 n262 GND GND nmos w=1u l=1u
M276 n259 N115 GND GND nmos w=1u l=1u
M277 n259 n262 net41 VDD pmos w=2u l=1u
M278 net41 N115 VDD VDD pmos w=2u l=1u
M279 n262 n213 GND GND nmos w=1u l=1u
M280 n262 n263 GND GND nmos w=1u l=1u
M281 n262 n213 net41 VDD pmos w=2u l=1u
M282 net41 n263 VDD VDD pmos w=2u l=1u
M283 n257 n239 n0 GND nmos w=1u l=1u
M284 n0 n264 GND GND nmos w=1u l=1u
M285 n257 n239 VDD VDD pmos w=2u l=1u
M286 n257 n264 VDD VDD pmos w=2u l=1u
M287 n239 n194 VDD VDD pmos w=2u l=1u
M288 n239 n194 GND GND nmos w=1u l=1u
M289 n264 n265 GND GND nmos w=1u l=1u
M290 n264 N53 GND GND nmos w=1u l=1u
M291 n264 n265 net41 VDD pmos w=2u l=1u
M292 net41 N53 VDD VDD pmos w=2u l=1u
M293 n265 n213 GND GND nmos w=1u l=1u
M294 n265 n193 GND GND nmos w=1u l=1u
M295 n265 n213 net41 VDD pmos w=2u l=1u
M296 net41 n193 VDD VDD pmos w=2u l=1u
M297 n255 n267 n0 GND nmos w=1u l=1u
M298 n0 n266 GND GND nmos w=1u l=1u
M299 n255 n267 VDD VDD pmos w=2u l=1u
M300 n255 n266 VDD VDD pmos w=2u l=1u
M301 n267 n269 n0 GND nmos w=1u l=1u
M302 n0 n268 GND GND nmos w=1u l=1u
M303 n267 n269 VDD VDD pmos w=2u l=1u
M304 n267 n268 VDD VDD pmos w=2u l=1u
M305 n269 n270 GND GND nmos w=1u l=1u
M306 n269 N14 GND GND nmos w=1u l=1u
M307 n269 n270 net41 VDD pmos w=2u l=1u
M308 net41 N14 VDD VDD pmos w=2u l=1u
M309 n268 n272 GND GND nmos w=1u l=1u
M310 n268 n271 GND GND nmos w=1u l=1u
M311 n268 n272 net41 VDD pmos w=2u l=1u
M312 net41 n271 VDD VDD pmos w=2u l=1u
M313 n271 n0 GND GND nmos w=1u l=1u
M314 net127 N8 GND GND nmos w=1u l=1u
M315 n0 N329 net127 GND nmos w=1u l=1u
M316 n0 N8 VDD VDD pmos w=2u l=1u
M317 n0 N329 VDD VDD pmos w=2u l=1u
M318 n271 n0 VDD VDD pmos w=2u l=1u
M319 n266 n274 GND GND nmos w=1u l=1u
M320 n266 n273 GND GND nmos w=1u l=1u
M321 n266 n274 net41 VDD pmos w=2u l=1u
M322 net41 n273 VDD VDD pmos w=2u l=1u
M323 n274 n275 GND GND nmos w=1u l=1u
M324 n274 n217 GND GND nmos w=1u l=1u
M325 n274 n275 net41 VDD pmos w=2u l=1u
M326 net41 n217 VDD VDD pmos w=2u l=1u
M327 n275 n220 n0 GND nmos w=1u l=1u
M328 n0 n276 GND GND nmos w=1u l=1u
M329 n275 n220 VDD VDD pmos w=2u l=1u
M330 n275 n276 VDD VDD pmos w=2u l=1u
M331 n220 N92 VDD VDD pmos w=2u l=1u
M332 n220 N92 GND GND nmos w=1u l=1u
M333 n276 n0 GND GND nmos w=1u l=1u
M334 n0 n213 GND GND nmos w=1u l=1u
M335 n0 n277 GND GND nmos w=1u l=1u
M336 n0 n277 n1 VDD pmos w=2u l=1u
M337 n276 n0 VDD VDD pmos w=2u l=1u
M338 n1 n213 VDD VDD pmos w=2u l=1u
M339 n273 n279 GND GND nmos w=1u l=1u
M340 n273 n278 GND GND nmos w=1u l=1u
M341 n273 n279 net41 VDD pmos w=2u l=1u
M342 net41 n278 VDD VDD pmos w=2u l=1u
M343 n279 n212 n0 GND nmos w=1u l=1u
M344 n0 n280 GND GND nmos w=1u l=1u
M345 n279 n212 VDD VDD pmos w=2u l=1u
M346 n279 n280 VDD VDD pmos w=2u l=1u
M347 n212 N105 VDD VDD pmos w=2u l=1u
M348 n212 N105 GND GND nmos w=1u l=1u
M349 n280 n281 n0 GND nmos w=1u l=1u
M350 n0 N329 GND GND nmos w=1u l=1u
M351 n280 n281 VDD VDD pmos w=2u l=1u
M352 n280 N329 VDD VDD pmos w=2u l=1u
M353 n253 n283 GND GND nmos w=1u l=1u
M354 n253 n282 GND GND nmos w=1u l=1u
M355 n253 n283 net41 VDD pmos w=2u l=1u
M356 net41 n282 VDD VDD pmos w=2u l=1u
M357 n283 n285 n0 GND nmos w=1u l=1u
M358 n0 n284 GND GND nmos w=1u l=1u
M359 n283 n285 VDD VDD pmos w=2u l=1u
M360 n283 n284 VDD VDD pmos w=2u l=1u
M361 n285 n287 n0 GND nmos w=1u l=1u
M362 n0 n286 GND GND nmos w=1u l=1u
M363 n285 n287 VDD VDD pmos w=2u l=1u
M364 n285 n286 VDD VDD pmos w=2u l=1u
M365 n287 n288 GND GND nmos w=1u l=1u
M366 n287 N27 GND GND nmos w=1u l=1u
M367 n287 n288 net41 VDD pmos w=2u l=1u
M368 net41 N27 VDD VDD pmos w=2u l=1u
M369 n288 n0 GND GND nmos w=1u l=1u
M370 net127 N329 GND GND nmos w=1u l=1u
M371 n0 n289 net127 GND nmos w=1u l=1u
M372 n0 N329 VDD VDD pmos w=2u l=1u
M373 n0 n289 VDD VDD pmos w=2u l=1u
M374 n288 n0 VDD VDD pmos w=2u l=1u
M375 n286 n291 GND GND nmos w=1u l=1u
M376 n286 n290 GND GND nmos w=1u l=1u
M377 n286 n291 net41 VDD pmos w=2u l=1u
M378 net41 n290 VDD VDD pmos w=2u l=1u
M379 n291 N17 VDD VDD pmos w=2u l=1u
M380 n291 N17 GND GND nmos w=1u l=1u
M381 n290 n293 GND GND nmos w=1u l=1u
M382 n290 n292 GND GND nmos w=1u l=1u
M383 n290 n293 net41 VDD pmos w=2u l=1u
M384 net41 n292 VDD VDD pmos w=2u l=1u
M385 n284 n295 n0 GND nmos w=1u l=1u
M386 n0 n294 GND GND nmos w=1u l=1u
M387 n284 n295 VDD VDD pmos w=2u l=1u
M388 n284 n294 VDD VDD pmos w=2u l=1u
M389 n295 n244 GND GND nmos w=1u l=1u
M390 n295 N40 GND GND nmos w=1u l=1u
M391 n295 n244 net41 VDD pmos w=2u l=1u
M392 net41 N40 VDD VDD pmos w=2u l=1u
M393 n294 n247 GND GND nmos w=1u l=1u
M394 n294 n296 GND GND nmos w=1u l=1u
M395 n294 n247 net41 VDD pmos w=2u l=1u
M396 net41 n296 VDD VDD pmos w=2u l=1u
M397 n296 n0 GND GND nmos w=1u l=1u
M398 net127 N329 GND GND nmos w=1u l=1u
M399 n0 n297 net127 GND nmos w=1u l=1u
M400 n0 N329 VDD VDD pmos w=2u l=1u
M401 n0 n297 VDD VDD pmos w=2u l=1u
M402 n296 n0 VDD VDD pmos w=2u l=1u
M403 n282 n299 n0 GND nmos w=1u l=1u
M404 n0 n298 GND GND nmos w=1u l=1u
M405 n282 n299 VDD VDD pmos w=2u l=1u
M406 n282 n298 VDD VDD pmos w=2u l=1u
M407 n299 n222 n0 GND nmos w=1u l=1u
M408 n0 n300 GND GND nmos w=1u l=1u
M409 n299 n222 VDD VDD pmos w=2u l=1u
M410 n299 n300 VDD VDD pmos w=2u l=1u
M411 n300 n301 GND GND nmos w=1u l=1u
M412 n300 N79 GND GND nmos w=1u l=1u
M413 n300 n301 net41 VDD pmos w=2u l=1u
M414 net41 N79 VDD VDD pmos w=2u l=1u
M415 n301 n213 GND GND nmos w=1u l=1u
M416 n301 n302 GND GND nmos w=1u l=1u
M417 n301 n213 net41 VDD pmos w=2u l=1u
M418 net41 n302 VDD VDD pmos w=2u l=1u
M419 n213 N329 VDD VDD pmos w=2u l=1u
M420 n213 N329 GND GND nmos w=1u l=1u
M421 n298 n234 n0 GND nmos w=1u l=1u
M422 n0 n303 GND GND nmos w=1u l=1u
M423 n298 n234 VDD VDD pmos w=2u l=1u
M424 n298 n303 VDD VDD pmos w=2u l=1u
M425 n303 n304 GND GND nmos w=1u l=1u
M426 n303 N66 GND GND nmos w=1u l=1u
M427 n303 n304 net41 VDD pmos w=2u l=1u
M428 net41 N66 VDD VDD pmos w=2u l=1u
M429 n304 n0 GND GND nmos w=1u l=1u
M430 net127 N329 GND GND nmos w=1u l=1u
M431 n0 n305 net127 GND nmos w=1u l=1u
M432 n0 N329 VDD VDD pmos w=2u l=1u
M433 n0 n305 VDD VDD pmos w=2u l=1u
M434 n304 n0 VDD VDD pmos w=2u l=1u
M435 N329 n307 n0 GND nmos w=1u l=1u
M436 n0 n306 GND GND nmos w=1u l=1u
M437 N329 n307 VDD VDD pmos w=2u l=1u
M438 N329 n306 VDD VDD pmos w=2u l=1u
M439 n307 n309 GND GND nmos w=1u l=1u
M440 n307 n308 GND GND nmos w=1u l=1u
M441 n307 n309 net41 VDD pmos w=2u l=1u
M442 net41 n308 VDD VDD pmos w=2u l=1u
M443 n309 n281 n0 GND nmos w=1u l=1u
M444 n0 n289 GND GND nmos w=1u l=1u
M445 n309 n281 VDD VDD pmos w=2u l=1u
M446 n309 n289 VDD VDD pmos w=2u l=1u
M447 n281 n214 n0 GND nmos w=1u l=1u
M448 n0 n208 GND GND nmos w=1u l=1u
M449 n281 n214 VDD VDD pmos w=2u l=1u
M450 n281 n208 VDD VDD pmos w=2u l=1u
M451 n214 N99 VDD VDD pmos w=2u l=1u
M452 n214 N99 GND GND nmos w=1u l=1u
M453 n208 n278 VDD VDD pmos w=2u l=1u
M454 n208 n278 GND GND nmos w=1u l=1u
M455 n278 n310 n0 GND nmos w=1u l=1u
M456 n0 N95 GND GND nmos w=1u l=1u
M457 n278 n310 VDD VDD pmos w=2u l=1u
M458 n278 N95 VDD VDD pmos w=2u l=1u
M459 n310 N223 n0 GND nmos w=1u l=1u
M460 n0 N89 GND GND nmos w=1u l=1u
M461 n310 N223 VDD VDD pmos w=2u l=1u
M462 n310 N89 VDD VDD pmos w=2u l=1u
M463 n289 n232 n0 GND nmos w=1u l=1u
M464 n0 n229 GND GND nmos w=1u l=1u
M465 n289 n232 VDD VDD pmos w=2u l=1u
M466 n289 n229 VDD VDD pmos w=2u l=1u
M467 n232 N21 VDD VDD pmos w=2u l=1u
M468 n232 N21 GND GND nmos w=1u l=1u
M469 n229 n0 GND GND nmos w=1u l=1u
M470 net127 n311 GND GND nmos w=1u l=1u
M471 n0 N17 net127 GND nmos w=1u l=1u
M472 n0 n311 VDD VDD pmos w=2u l=1u
M473 n0 N17 VDD VDD pmos w=2u l=1u
M474 n229 n0 VDD VDD pmos w=2u l=1u
M475 n311 N223 n0 GND nmos w=1u l=1u
M476 n0 N11 GND GND nmos w=1u l=1u
M477 n311 N223 VDD VDD pmos w=2u l=1u
M478 n311 N11 VDD VDD pmos w=2u l=1u
M479 n308 n313 n0 GND nmos w=1u l=1u
M480 n0 n312 GND GND nmos w=1u l=1u
M481 n308 n313 VDD VDD pmos w=2u l=1u
M482 n308 n312 VDD VDD pmos w=2u l=1u
M483 n313 n263 VDD VDD pmos w=2u l=1u
M484 n313 n263 GND GND nmos w=1u l=1u
M485 n263 n261 GND GND nmos w=1u l=1u
M486 n263 N112 GND GND nmos w=1u l=1u
M487 n263 n261 net41 VDD pmos w=2u l=1u
M488 net41 N112 VDD VDD pmos w=2u l=1u
M489 n261 n314 n0 GND nmos w=1u l=1u
M490 n0 N108 GND GND nmos w=1u l=1u
M491 n261 n314 VDD VDD pmos w=2u l=1u
M492 n261 N108 VDD VDD pmos w=2u l=1u
M493 n314 N223 n0 GND nmos w=1u l=1u
M494 n0 N102 GND GND nmos w=1u l=1u
M495 n314 N223 VDD VDD pmos w=2u l=1u
M496 n314 N102 VDD VDD pmos w=2u l=1u
M497 n312 n302 GND GND nmos w=1u l=1u
M498 n312 n277 GND GND nmos w=1u l=1u
M499 n312 n302 net41 VDD pmos w=2u l=1u
M500 net41 n277 VDD VDD pmos w=2u l=1u
M501 n302 n0 GND GND nmos w=1u l=1u
M502 net127 n225 GND GND nmos w=1u l=1u
M503 n0 n222 net127 GND nmos w=1u l=1u
M504 n0 n225 VDD VDD pmos w=2u l=1u
M505 n0 n222 VDD VDD pmos w=2u l=1u
M506 n302 n0 VDD VDD pmos w=2u l=1u
M507 n225 N73 VDD VDD pmos w=2u l=1u
M508 n225 N73 GND GND nmos w=1u l=1u
M509 n222 n0 GND GND nmos w=1u l=1u
M510 net127 n315 GND GND nmos w=1u l=1u
M511 n0 N69 net127 GND nmos w=1u l=1u
M512 n0 n315 VDD VDD pmos w=2u l=1u
M513 n0 N69 VDD VDD pmos w=2u l=1u
M514 n222 n0 VDD VDD pmos w=2u l=1u
M515 n315 N223 n0 GND nmos w=1u l=1u
M516 n0 N63 GND GND nmos w=1u l=1u
M517 n315 N223 VDD VDD pmos w=2u l=1u
M518 n315 N63 VDD VDD pmos w=2u l=1u
M519 n277 N86 GND GND nmos w=1u l=1u
M520 n277 n217 GND GND nmos w=1u l=1u
M521 n277 N86 net41 VDD pmos w=2u l=1u
M522 net41 n217 VDD VDD pmos w=2u l=1u
M523 n217 n316 n0 GND nmos w=1u l=1u
M524 n0 N82 GND GND nmos w=1u l=1u
M525 n217 n316 VDD VDD pmos w=2u l=1u
M526 n217 N82 VDD VDD pmos w=2u l=1u
M527 n316 N223 n0 GND nmos w=1u l=1u
M528 n0 N76 GND GND nmos w=1u l=1u
M529 n316 N223 VDD VDD pmos w=2u l=1u
M530 n316 N76 VDD VDD pmos w=2u l=1u
M531 n306 n318 GND GND nmos w=1u l=1u
M532 n306 n317 GND GND nmos w=1u l=1u
M533 n306 n318 net41 VDD pmos w=2u l=1u
M534 net41 n317 VDD VDD pmos w=2u l=1u
M535 n318 n320 n0 GND nmos w=1u l=1u
M536 n0 n319 GND GND nmos w=1u l=1u
M537 n318 n320 VDD VDD pmos w=2u l=1u
M538 n318 n319 VDD VDD pmos w=2u l=1u
M539 n320 n193 VDD VDD pmos w=2u l=1u
M540 n320 n193 GND GND nmos w=1u l=1u
M541 n193 N47 GND GND nmos w=1u l=1u
M542 n193 n194 GND GND nmos w=1u l=1u
M543 n193 N47 net41 VDD pmos w=2u l=1u
M544 net41 n194 VDD VDD pmos w=2u l=1u
M545 n194 n321 n0 GND nmos w=1u l=1u
M546 n0 N43 GND GND nmos w=1u l=1u
M547 n194 n321 VDD VDD pmos w=2u l=1u
M548 n194 N43 VDD VDD pmos w=2u l=1u
M549 n321 N223 n0 GND nmos w=1u l=1u
M550 n0 N37 GND GND nmos w=1u l=1u
M551 n321 N223 VDD VDD pmos w=2u l=1u
M552 n321 N37 VDD VDD pmos w=2u l=1u
M553 n319 N4 n0 GND nmos w=1u l=1u
M554 n0 n322 GND GND nmos w=1u l=1u
M555 n319 N4 VDD VDD pmos w=2u l=1u
M556 n319 n322 VDD VDD pmos w=2u l=1u
M557 n322 n270 GND GND nmos w=1u l=1u
M558 n322 N8 GND GND nmos w=1u l=1u
M559 n322 n270 net41 VDD pmos w=2u l=1u
M560 net41 N8 VDD VDD pmos w=2u l=1u
M561 n270 n252 VDD VDD pmos w=2u l=1u
M562 n270 n252 GND GND nmos w=1u l=1u
M563 n252 N223 n0 GND nmos w=1u l=1u
M564 n0 N1 GND GND nmos w=1u l=1u
M565 n252 N223 VDD VDD pmos w=2u l=1u
M566 n252 N1 VDD VDD pmos w=2u l=1u
M567 n317 n297 n0 GND nmos w=1u l=1u
M568 n0 n305 GND GND nmos w=1u l=1u
M569 n317 n297 VDD VDD pmos w=2u l=1u
M570 n317 n305 VDD VDD pmos w=2u l=1u
M571 n297 N30 n0 GND nmos w=1u l=1u
M572 n0 n323 GND GND nmos w=1u l=1u
M573 n297 N30 VDD VDD pmos w=2u l=1u
M574 n297 n323 VDD VDD pmos w=2u l=1u
M575 n323 n244 GND GND nmos w=1u l=1u
M576 n323 N34 GND GND nmos w=1u l=1u
M577 n323 n244 net41 VDD pmos w=2u l=1u
M578 net41 N34 VDD VDD pmos w=2u l=1u
M579 n244 n324 GND GND nmos w=1u l=1u
M580 n244 n292 GND GND nmos w=1u l=1u
M581 n244 n324 net41 VDD pmos w=2u l=1u
M582 net41 n292 VDD VDD pmos w=2u l=1u
M583 n292 N223 VDD VDD pmos w=2u l=1u
M584 n292 N223 GND GND nmos w=1u l=1u
M585 n305 n237 n0 GND nmos w=1u l=1u
M586 n0 n234 GND GND nmos w=1u l=1u
M587 n305 n237 VDD VDD pmos w=2u l=1u
M588 n305 n234 VDD VDD pmos w=2u l=1u
M589 n237 N60 VDD VDD pmos w=2u l=1u
M590 n237 N60 GND GND nmos w=1u l=1u
M591 n234 n0 GND GND nmos w=1u l=1u
M592 net127 n325 GND GND nmos w=1u l=1u
M593 n0 N56 net127 GND nmos w=1u l=1u
M594 n0 n325 VDD VDD pmos w=2u l=1u
M595 n0 N56 VDD VDD pmos w=2u l=1u
M596 n234 n0 VDD VDD pmos w=2u l=1u
M597 n325 N223 n0 GND nmos w=1u l=1u
M598 n0 N50 GND GND nmos w=1u l=1u
M599 n325 N223 VDD VDD pmos w=2u l=1u
M600 n325 N50 VDD VDD pmos w=2u l=1u
M601 N223 n327 n0 GND nmos w=1u l=1u
M602 n0 n326 GND GND nmos w=1u l=1u
M603 N223 n327 VDD VDD pmos w=2u l=1u
M604 N223 n326 VDD VDD pmos w=2u l=1u
M605 n327 n329 GND GND nmos w=1u l=1u
M606 n327 n328 GND GND nmos w=1u l=1u
M607 n327 n329 net41 VDD pmos w=2u l=1u
M608 net41 n328 VDD VDD pmos w=2u l=1u
M609 n329 n331 n0 GND nmos w=1u l=1u
M610 n0 n330 GND GND nmos w=1u l=1u
M611 n329 n331 VDD VDD pmos w=2u l=1u
M612 n329 n330 VDD VDD pmos w=2u l=1u
M613 n331 n293 n0 GND nmos w=1u l=1u
M614 n0 N17 GND GND nmos w=1u l=1u
M615 n331 n293 VDD VDD pmos w=2u l=1u
M616 n331 N17 VDD VDD pmos w=2u l=1u
M617 n293 N11 VDD VDD pmos w=2u l=1u
M618 n293 N11 GND GND nmos w=1u l=1u
M619 n330 n332 n0 GND nmos w=1u l=1u
M620 n0 N43 GND GND nmos w=1u l=1u
M621 n330 n332 VDD VDD pmos w=2u l=1u
M622 n330 N43 VDD VDD pmos w=2u l=1u
M623 n332 N37 VDD VDD pmos w=2u l=1u
M624 n332 N37 GND GND nmos w=1u l=1u
M625 n328 n334 n0 GND nmos w=1u l=1u
M626 n0 n333 GND GND nmos w=1u l=1u
M627 n328 n334 VDD VDD pmos w=2u l=1u
M628 n328 n333 VDD VDD pmos w=2u l=1u
M629 n334 n335 n0 GND nmos w=1u l=1u
M630 n0 N108 GND GND nmos w=1u l=1u
M631 n334 n335 VDD VDD pmos w=2u l=1u
M632 n334 N108 VDD VDD pmos w=2u l=1u
M633 n335 N102 VDD VDD pmos w=2u l=1u
M634 n335 N102 GND GND nmos w=1u l=1u
M635 n333 n336 GND GND nmos w=1u l=1u
M636 n333 n324 GND GND nmos w=1u l=1u
M637 n333 n336 net41 VDD pmos w=2u l=1u
M638 net41 n324 VDD VDD pmos w=2u l=1u
M639 n336 n272 GND GND nmos w=1u l=1u
M640 n336 N1 GND GND nmos w=1u l=1u
M641 n336 n272 net41 VDD pmos w=2u l=1u
M642 net41 N1 VDD VDD pmos w=2u l=1u
M643 n272 N4 VDD VDD pmos w=2u l=1u
M644 n272 N4 GND GND nmos w=1u l=1u
M645 n324 n247 GND GND nmos w=1u l=1u
M646 n324 N24 GND GND nmos w=1u l=1u
M647 n324 n247 net41 VDD pmos w=2u l=1u
M648 net41 N24 VDD VDD pmos w=2u l=1u
M649 n247 N30 VDD VDD pmos w=2u l=1u
M650 n247 N30 GND GND nmos w=1u l=1u
M651 n326 n338 GND GND nmos w=1u l=1u
M652 n326 n337 GND GND nmos w=1u l=1u
M653 n326 n338 net41 VDD pmos w=2u l=1u
M654 net41 n337 VDD VDD pmos w=2u l=1u
M655 n338 n340 n0 GND nmos w=1u l=1u
M656 n0 n339 GND GND nmos w=1u l=1u
M657 n338 n340 VDD VDD pmos w=2u l=1u
M658 n338 n339 VDD VDD pmos w=2u l=1u
M659 n340 n341 n0 GND nmos w=1u l=1u
M660 n0 N82 GND GND nmos w=1u l=1u
M661 n340 n341 VDD VDD pmos w=2u l=1u
M662 n340 N82 VDD VDD pmos w=2u l=1u
M663 n341 N76 VDD VDD pmos w=2u l=1u
M664 n341 N76 GND GND nmos w=1u l=1u
M665 n339 n342 n0 GND nmos w=1u l=1u
M666 n0 N95 GND GND nmos w=1u l=1u
M667 n339 n342 VDD VDD pmos w=2u l=1u
M668 n339 N95 VDD VDD pmos w=2u l=1u
M669 n342 N89 VDD VDD pmos w=2u l=1u
M670 n342 N89 GND GND nmos w=1u l=1u
M671 n337 n344 n0 GND nmos w=1u l=1u
M672 n0 n343 GND GND nmos w=1u l=1u
M673 n337 n344 VDD VDD pmos w=2u l=1u
M674 n337 n343 VDD VDD pmos w=2u l=1u
M675 n344 n345 n0 GND nmos w=1u l=1u
M676 n0 N56 GND GND nmos w=1u l=1u
M677 n344 n345 VDD VDD pmos w=2u l=1u
M678 n344 N56 VDD VDD pmos w=2u l=1u
M679 n345 N50 VDD VDD pmos w=2u l=1u
M680 n345 N50 GND GND nmos w=1u l=1u
M681 n343 n346 n0 GND nmos w=1u l=1u
M682 n0 N69 GND GND nmos w=1u l=1u
M683 n343 n346 VDD VDD pmos w=2u l=1u
M684 n343 N69 VDD VDD pmos w=2u l=1u
M685 n346 N63 VDD VDD pmos w=2u l=1u
M686 n346 N63 GND GND nmos w=1u l=1u
.ENDS


