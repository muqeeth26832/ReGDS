.SUBCKT c6288 N1 N18 N35 N52 N69 N86 N103 N120 N137 N154 N171 N188 N205 N222 N239 N256 N273 N290 N307 N324 N341 N358 N375 N392 N409 N426 N443 N460 N477 N494 N511 N528 N545 N1581 N1901 N2223 N2548 N2877 N3211 N3552 N3895 N4241 N4591 N4946 N5308 N5672 N5971 N6123 N6150 N6160 N6170 N6180 N6190 N6200 N6210 N6220 N6230 N6240 N6250 N6260 N6270 N6280 N6287 N6288 VDD VSS 
M1 N6288 n2200 net1 VSS nmos w=1u l=1u
M2 net1 n2199 VSS VSS nmos w=1u l=1u
M3 N6288 n2200 VDD VDD pmos w=2u l=1u
M4 N6288 n2199 VDD VDD pmos w=2u l=1u
M5 n2200 n2202 net2 VSS nmos w=1u l=1u
M6 net2 n2201 VSS VSS nmos w=1u l=1u
M7 n2200 n2202 VDD VDD pmos w=2u l=1u
M8 n2200 n2201 VDD VDD pmos w=2u l=1u
M9 n2201 net3 VSS VSS nmos w=1u l=1u
M10 net4 n2204 VSS VSS nmos w=1u l=1u
M11 net3 n2203 net4 VSS nmos w=1u l=1u
M12 net3 n2204 VDD VDD pmos w=2u l=1u
M13 net3 n2203 VDD VDD pmos w=2u l=1u
M14 n2201 net3 VDD VDD pmos w=2u l=1u
M15 N6287 n2206 VSS VSS nmos w=1u l=1u
M16 N6287 n2205 VSS VSS nmos w=1u l=1u
M17 N6287 n2206 net5 VDD pmos w=2u l=1u
M18 net5 n2205 VDD VDD pmos w=2u l=1u
M19 n2206 n2199 net6 VSS nmos w=1u l=1u
M20 net6 N256 VSS VSS nmos w=1u l=1u
M21 n2206 n2199 VDD VDD pmos w=2u l=1u
M22 n2206 N256 VDD VDD pmos w=2u l=1u
M23 n2199 n2208 net7 VSS nmos w=1u l=1u
M24 net7 n2207 VSS VSS nmos w=1u l=1u
M25 n2199 n2208 VDD VDD pmos w=2u l=1u
M26 n2199 n2207 VDD VDD pmos w=2u l=1u
M27 n2208 n2203 net8 VSS nmos w=1u l=1u
M28 net8 n2204 VSS VSS nmos w=1u l=1u
M29 n2208 n2203 VDD VDD pmos w=2u l=1u
M30 n2208 n2204 VDD VDD pmos w=2u l=1u
M31 n2207 n2202 VDD VDD pmos w=2u l=1u
M32 n2207 n2202 VSS VSS nmos w=1u l=1u
M33 net9 n2210 VSS VSS nmos w=1u l=1u
M34 net10 n2209 VSS VSS nmos w=1u l=1u
M35 n2202 net11 VSS VSS nmos w=1u l=1u
M36 net11 n2210 net12 VSS nmos w=1u l=1u
M37 net11 net9 net10 VSS nmos w=1u l=1u
M38 net12 net10 VSS VSS nmos w=1u l=1u
M39 net11 net9 net13 VDD pmos w=2u l=1u
M40 net9 n2210 VDD VDD pmos w=2u l=1u
M41 net10 n2210 net11 VDD pmos w=2u l=1u
M42 net10 n2209 VDD VDD pmos w=2u l=1u
M43 n2202 net11 VDD VDD pmos w=2u l=1u
M44 net13 net10 VDD VDD pmos w=2u l=1u
M45 n2210 net14 VSS VSS nmos w=1u l=1u
M46 net15 n2212 VSS VSS nmos w=1u l=1u
M47 net14 n2211 net15 VSS nmos w=1u l=1u
M48 net14 n2212 VDD VDD pmos w=2u l=1u
M49 net14 n2211 VDD VDD pmos w=2u l=1u
M50 n2210 net14 VDD VDD pmos w=2u l=1u
M51 n2209 N256 net16 VSS nmos w=1u l=1u
M52 net16 N528 VSS VSS nmos w=1u l=1u
M53 n2209 N256 VDD VDD pmos w=2u l=1u
M54 n2209 N528 VDD VDD pmos w=2u l=1u
M55 N6280 n2213 net17 VSS nmos w=1u l=1u
M56 net17 n2204 VSS VSS nmos w=1u l=1u
M57 N6280 n2213 VDD VDD pmos w=2u l=1u
M58 N6280 n2204 VDD VDD pmos w=2u l=1u
M59 n2213 n2215 net18 VSS nmos w=1u l=1u
M60 net18 n2214 VSS VSS nmos w=1u l=1u
M61 n2213 n2215 VDD VDD pmos w=2u l=1u
M62 n2213 n2214 VDD VDD pmos w=2u l=1u
M63 n2214 n2217 VSS VSS nmos w=1u l=1u
M64 n2214 n2216 VSS VSS nmos w=1u l=1u
M65 n2214 n2217 net19 VDD pmos w=2u l=1u
M66 net19 n2216 VDD VDD pmos w=2u l=1u
M67 n2216 n2218 VDD VDD pmos w=2u l=1u
M68 n2216 n2218 VSS VSS nmos w=1u l=1u
M69 n2204 n2219 net20 VSS nmos w=1u l=1u
M70 net20 n2217 VSS VSS nmos w=1u l=1u
M71 n2204 n2219 VDD VDD pmos w=2u l=1u
M72 n2204 n2217 VDD VDD pmos w=2u l=1u
M73 n2219 n2218 net21 VSS nmos w=1u l=1u
M74 net21 n2215 VSS VSS nmos w=1u l=1u
M75 n2219 n2218 VDD VDD pmos w=2u l=1u
M76 n2219 n2215 VDD VDD pmos w=2u l=1u
M77 n2217 net22 VSS VSS nmos w=1u l=1u
M78 net23 n2220 VSS VSS nmos w=1u l=1u
M79 net22 n2203 net23 VSS nmos w=1u l=1u
M80 net22 n2220 VDD VDD pmos w=2u l=1u
M81 net22 n2203 VDD VDD pmos w=2u l=1u
M82 n2217 net22 VDD VDD pmos w=2u l=1u
M83 n2220 n2222 net24 VSS nmos w=1u l=1u
M84 net24 n2221 VSS VSS nmos w=1u l=1u
M85 n2220 n2222 VDD VDD pmos w=2u l=1u
M86 n2220 n2221 VDD VDD pmos w=2u l=1u
M87 n2203 net25 VSS VSS nmos w=1u l=1u
M88 net25 n2222 VSS VSS nmos w=1u l=1u
M89 net25 n2221 VSS VSS nmos w=1u l=1u
M90 net25 n2221 net26 VDD pmos w=2u l=1u
M91 n2203 net25 VDD VDD pmos w=2u l=1u
M92 net26 n2222 VDD VDD pmos w=2u l=1u
M93 n2221 net27 VSS VSS nmos w=1u l=1u
M94 net28 n2224 VSS VSS nmos w=1u l=1u
M95 net27 n2223 net28 VSS nmos w=1u l=1u
M96 net27 n2224 VDD VDD pmos w=2u l=1u
M97 net27 n2223 VDD VDD pmos w=2u l=1u
M98 n2221 net27 VDD VDD pmos w=2u l=1u
M99 n2222 n2225 net29 VSS nmos w=1u l=1u
M100 net29 n2212 VSS VSS nmos w=1u l=1u
M101 n2222 n2225 VDD VDD pmos w=2u l=1u
M102 n2222 n2212 VDD VDD pmos w=2u l=1u
M103 n2225 N528 net30 VSS nmos w=1u l=1u
M104 net30 n2226 VSS VSS nmos w=1u l=1u
M105 n2225 N528 VDD VDD pmos w=2u l=1u
M106 n2225 n2226 VDD VDD pmos w=2u l=1u
M107 n2226 n2228 VSS VSS nmos w=1u l=1u
M108 n2226 n2227 VSS VSS nmos w=1u l=1u
M109 n2226 n2228 net31 VDD pmos w=2u l=1u
M110 net31 n2227 VDD VDD pmos w=2u l=1u
M111 n2212 n2229 net32 VSS nmos w=1u l=1u
M112 net32 n2227 VSS VSS nmos w=1u l=1u
M113 n2212 n2229 VDD VDD pmos w=2u l=1u
M114 n2212 n2227 VDD VDD pmos w=2u l=1u
M115 n2229 N239 net33 VSS nmos w=1u l=1u
M116 net33 N528 VSS VSS nmos w=1u l=1u
M117 n2229 N239 VDD VDD pmos w=2u l=1u
M118 n2229 N528 VDD VDD pmos w=2u l=1u
M119 n2227 net34 VSS VSS nmos w=1u l=1u
M120 net35 n2230 VSS VSS nmos w=1u l=1u
M121 net34 n2211 net35 VSS nmos w=1u l=1u
M122 net34 n2230 VDD VDD pmos w=2u l=1u
M123 net34 n2211 VDD VDD pmos w=2u l=1u
M124 n2227 net34 VDD VDD pmos w=2u l=1u
M125 n2230 net36 VSS VSS nmos w=1u l=1u
M126 net36 n2231 VSS VSS nmos w=1u l=1u
M127 net36 n2232 VSS VSS nmos w=1u l=1u
M128 net36 n2232 net37 VDD pmos w=2u l=1u
M129 n2230 net36 VDD VDD pmos w=2u l=1u
M130 net37 n2231 VDD VDD pmos w=2u l=1u
M131 n2211 n2233 net38 VSS nmos w=1u l=1u
M132 net38 n2231 VSS VSS nmos w=1u l=1u
M133 n2211 n2233 VDD VDD pmos w=2u l=1u
M134 n2211 n2231 VDD VDD pmos w=2u l=1u
M135 n2233 N511 net39 VSS nmos w=1u l=1u
M136 net39 N256 VSS VSS nmos w=1u l=1u
M137 n2233 N511 VDD VDD pmos w=2u l=1u
M138 n2233 N256 VDD VDD pmos w=2u l=1u
M139 n2231 n2235 net40 VSS nmos w=1u l=1u
M140 net40 n2234 VSS VSS nmos w=1u l=1u
M141 n2231 n2235 VDD VDD pmos w=2u l=1u
M142 n2231 n2234 VDD VDD pmos w=2u l=1u
M143 n2234 n2237 net41 VSS nmos w=1u l=1u
M144 net41 n2236 VSS VSS nmos w=1u l=1u
M145 n2234 n2237 VDD VDD pmos w=2u l=1u
M146 n2234 n2236 VDD VDD pmos w=2u l=1u
M147 n2237 N256 net42 VSS nmos w=1u l=1u
M148 net42 N494 VSS VSS nmos w=1u l=1u
M149 n2237 N256 VDD VDD pmos w=2u l=1u
M150 n2237 N494 VDD VDD pmos w=2u l=1u
M151 N6270 n2238 net43 VSS nmos w=1u l=1u
M152 net43 n2218 VSS VSS nmos w=1u l=1u
M153 N6270 n2238 VDD VDD pmos w=2u l=1u
M154 N6270 n2218 VDD VDD pmos w=2u l=1u
M155 n2238 n2240 net44 VSS nmos w=1u l=1u
M156 net44 n2239 VSS VSS nmos w=1u l=1u
M157 n2238 n2240 VDD VDD pmos w=2u l=1u
M158 n2238 n2239 VDD VDD pmos w=2u l=1u
M159 n2240 n2241 net45 VSS nmos w=1u l=1u
M160 net45 n2215 VSS VSS nmos w=1u l=1u
M161 n2240 n2241 VDD VDD pmos w=2u l=1u
M162 n2240 n2215 VDD VDD pmos w=2u l=1u
M163 n2241 n2243 net46 VSS nmos w=1u l=1u
M164 net46 n2242 VSS VSS nmos w=1u l=1u
M165 n2241 n2243 VDD VDD pmos w=2u l=1u
M166 n2241 n2242 VDD VDD pmos w=2u l=1u
M167 n2215 net47 VSS VSS nmos w=1u l=1u
M168 net47 n2243 VSS VSS nmos w=1u l=1u
M169 net47 n2242 VSS VSS nmos w=1u l=1u
M170 net47 n2242 net48 VDD pmos w=2u l=1u
M171 n2215 net47 VDD VDD pmos w=2u l=1u
M172 net48 n2243 VDD VDD pmos w=2u l=1u
M173 n2239 n2244 VDD VDD pmos w=2u l=1u
M174 n2239 n2244 VSS VSS nmos w=1u l=1u
M175 n2218 n2244 net49 VSS nmos w=1u l=1u
M176 net49 n2245 VSS VSS nmos w=1u l=1u
M177 n2218 n2244 VDD VDD pmos w=2u l=1u
M178 n2218 n2245 VDD VDD pmos w=2u l=1u
M179 n2244 n2247 net50 VSS nmos w=1u l=1u
M180 net50 n2246 VSS VSS nmos w=1u l=1u
M181 n2244 n2247 VDD VDD pmos w=2u l=1u
M182 n2244 n2246 VDD VDD pmos w=2u l=1u
M183 n2246 n2249 net51 VSS nmos w=1u l=1u
M184 net51 n2248 VSS VSS nmos w=1u l=1u
M185 n2246 n2249 VDD VDD pmos w=2u l=1u
M186 n2246 n2248 VDD VDD pmos w=2u l=1u
M187 net52 n2243 VSS VSS nmos w=1u l=1u
M188 net53 n2242 VSS VSS nmos w=1u l=1u
M189 n2245 net54 VSS VSS nmos w=1u l=1u
M190 net54 n2243 net55 VSS nmos w=1u l=1u
M191 net54 net52 net53 VSS nmos w=1u l=1u
M192 net55 net53 VSS VSS nmos w=1u l=1u
M193 net54 net52 net56 VDD pmos w=2u l=1u
M194 net52 n2243 VDD VDD pmos w=2u l=1u
M195 net53 n2243 net54 VDD pmos w=2u l=1u
M196 net53 n2242 VDD VDD pmos w=2u l=1u
M197 n2245 net54 VDD VDD pmos w=2u l=1u
M198 net56 net53 VDD VDD pmos w=2u l=1u
M199 n2243 n2250 net57 VSS nmos w=1u l=1u
M200 net57 n2224 VSS VSS nmos w=1u l=1u
M201 n2243 n2250 VDD VDD pmos w=2u l=1u
M202 n2243 n2224 VDD VDD pmos w=2u l=1u
M203 n2250 N222 net58 VSS nmos w=1u l=1u
M204 net58 n2251 VSS VSS nmos w=1u l=1u
M205 n2250 N222 VDD VDD pmos w=2u l=1u
M206 n2250 n2251 VDD VDD pmos w=2u l=1u
M207 n2251 n2205 VSS VSS nmos w=1u l=1u
M208 n2251 n2252 VSS VSS nmos w=1u l=1u
M209 n2251 n2205 net59 VDD pmos w=2u l=1u
M210 net59 n2252 VDD VDD pmos w=2u l=1u
M211 n2224 n2253 net60 VSS nmos w=1u l=1u
M212 net60 n2252 VSS VSS nmos w=1u l=1u
M213 n2224 n2253 VDD VDD pmos w=2u l=1u
M214 n2224 n2252 VDD VDD pmos w=2u l=1u
M215 n2253 N528 net61 VSS nmos w=1u l=1u
M216 net61 N222 VSS VSS nmos w=1u l=1u
M217 n2253 N528 VDD VDD pmos w=2u l=1u
M218 n2253 N222 VDD VDD pmos w=2u l=1u
M219 n2252 net62 VSS VSS nmos w=1u l=1u
M220 net63 n2223 VSS VSS nmos w=1u l=1u
M221 net62 n2254 net63 VSS nmos w=1u l=1u
M222 net62 n2223 VDD VDD pmos w=2u l=1u
M223 net62 n2254 VDD VDD pmos w=2u l=1u
M224 n2252 net62 VDD VDD pmos w=2u l=1u
M225 n2223 n2256 net64 VSS nmos w=1u l=1u
M226 net64 n2255 VSS VSS nmos w=1u l=1u
M227 n2223 n2256 VDD VDD pmos w=2u l=1u
M228 n2223 n2255 VDD VDD pmos w=2u l=1u
M229 n2256 n2258 net65 VSS nmos w=1u l=1u
M230 net65 n2257 VSS VSS nmos w=1u l=1u
M231 n2256 n2258 VDD VDD pmos w=2u l=1u
M232 n2256 n2257 VDD VDD pmos w=2u l=1u
M233 n2254 n2257 net66 VSS nmos w=1u l=1u
M234 net66 n2259 VSS VSS nmos w=1u l=1u
M235 n2254 n2257 VDD VDD pmos w=2u l=1u
M236 n2254 n2259 VDD VDD pmos w=2u l=1u
M237 n2257 n2261 net67 VSS nmos w=1u l=1u
M238 net67 n2260 VSS VSS nmos w=1u l=1u
M239 n2257 n2261 VDD VDD pmos w=2u l=1u
M240 n2257 n2260 VDD VDD pmos w=2u l=1u
M241 n2259 n2255 VSS VSS nmos w=1u l=1u
M242 n2259 n2262 VSS VSS nmos w=1u l=1u
M243 n2259 n2255 net68 VDD pmos w=2u l=1u
M244 net68 n2262 VDD VDD pmos w=2u l=1u
M245 n2255 net69 VSS VSS nmos w=1u l=1u
M246 net70 n2263 VSS VSS nmos w=1u l=1u
M247 net69 n2235 net70 VSS nmos w=1u l=1u
M248 net69 n2263 VDD VDD pmos w=2u l=1u
M249 net69 n2235 VDD VDD pmos w=2u l=1u
M250 n2255 net69 VDD VDD pmos w=2u l=1u
M251 n2263 N511 net71 VSS nmos w=1u l=1u
M252 net71 n2264 VSS VSS nmos w=1u l=1u
M253 n2263 N511 VDD VDD pmos w=2u l=1u
M254 n2263 n2264 VDD VDD pmos w=2u l=1u
M255 n2264 n2266 VSS VSS nmos w=1u l=1u
M256 n2264 n2265 VSS VSS nmos w=1u l=1u
M257 n2264 n2266 net72 VDD pmos w=2u l=1u
M258 net72 n2265 VDD VDD pmos w=2u l=1u
M259 n2266 n2268 VSS VSS nmos w=1u l=1u
M260 n2266 n2267 VSS VSS nmos w=1u l=1u
M261 n2266 n2268 net73 VDD pmos w=2u l=1u
M262 net73 n2267 VDD VDD pmos w=2u l=1u
M263 n2268 n2270 net74 VSS nmos w=1u l=1u
M264 net74 n2269 VSS VSS nmos w=1u l=1u
M265 n2268 n2270 VDD VDD pmos w=2u l=1u
M266 n2268 n2269 VDD VDD pmos w=2u l=1u
M267 n2269 n2271 net75 VSS nmos w=1u l=1u
M268 net75 N239 VSS VSS nmos w=1u l=1u
M269 n2269 n2271 VDD VDD pmos w=2u l=1u
M270 n2269 N239 VDD VDD pmos w=2u l=1u
M271 n2265 n2236 VSS VSS nmos w=1u l=1u
M272 n2265 N494 VSS VSS nmos w=1u l=1u
M273 n2265 n2236 net76 VDD pmos w=2u l=1u
M274 net76 N494 VDD VDD pmos w=2u l=1u
M275 n2235 n2273 net77 VSS nmos w=1u l=1u
M276 net77 n2272 VSS VSS nmos w=1u l=1u
M277 n2235 n2273 VDD VDD pmos w=2u l=1u
M278 n2235 n2272 VDD VDD pmos w=2u l=1u
M279 n2273 N239 net78 VSS nmos w=1u l=1u
M280 net78 N511 VSS VSS nmos w=1u l=1u
M281 n2273 N239 VDD VDD pmos w=2u l=1u
M282 n2273 N511 VDD VDD pmos w=2u l=1u
M283 net79 n2274 VSS VSS nmos w=1u l=1u
M284 net80 n2267 VSS VSS nmos w=1u l=1u
M285 n2272 net81 VSS VSS nmos w=1u l=1u
M286 net81 n2274 net82 VSS nmos w=1u l=1u
M287 net81 net79 net80 VSS nmos w=1u l=1u
M288 net82 net80 VSS VSS nmos w=1u l=1u
M289 net81 net79 net83 VDD pmos w=2u l=1u
M290 net79 n2274 VDD VDD pmos w=2u l=1u
M291 net80 n2274 net81 VDD pmos w=2u l=1u
M292 net80 n2267 VDD VDD pmos w=2u l=1u
M293 n2272 net81 VDD VDD pmos w=2u l=1u
M294 net83 net80 VDD VDD pmos w=2u l=1u
M295 n2274 n2271 VSS VSS nmos w=1u l=1u
M296 n2274 n2275 VSS VSS nmos w=1u l=1u
M297 n2274 n2271 net84 VDD pmos w=2u l=1u
M298 net84 n2275 VDD VDD pmos w=2u l=1u
M299 n2267 n2236 VDD VDD pmos w=2u l=1u
M300 n2267 n2236 VSS VSS nmos w=1u l=1u
M301 n2236 n2277 net85 VSS nmos w=1u l=1u
M302 net85 n2276 VSS VSS nmos w=1u l=1u
M303 n2236 n2277 VDD VDD pmos w=2u l=1u
M304 n2236 n2276 VDD VDD pmos w=2u l=1u
M305 n2277 n2279 net86 VSS nmos w=1u l=1u
M306 net86 n2278 VSS VSS nmos w=1u l=1u
M307 n2277 n2279 VDD VDD pmos w=2u l=1u
M308 n2277 n2278 VDD VDD pmos w=2u l=1u
M309 n2262 n2258 VDD VDD pmos w=2u l=1u
M310 n2262 n2258 VSS VSS nmos w=1u l=1u
M311 n2242 net87 VSS VSS nmos w=1u l=1u
M312 net88 n2281 VSS VSS nmos w=1u l=1u
M313 net87 n2280 net88 VSS nmos w=1u l=1u
M314 net87 n2281 VDD VDD pmos w=2u l=1u
M315 net87 n2280 VDD VDD pmos w=2u l=1u
M316 n2242 net87 VDD VDD pmos w=2u l=1u
M317 n2280 n2283 net89 VSS nmos w=1u l=1u
M318 net89 n2282 VSS VSS nmos w=1u l=1u
M319 n2280 n2283 VDD VDD pmos w=2u l=1u
M320 n2280 n2282 VDD VDD pmos w=2u l=1u
M321 N6260 n2284 net90 VSS nmos w=1u l=1u
M322 net90 n2247 VSS VSS nmos w=1u l=1u
M323 N6260 n2284 VDD VDD pmos w=2u l=1u
M324 N6260 n2247 VDD VDD pmos w=2u l=1u
M325 n2284 net91 VSS VSS nmos w=1u l=1u
M326 net91 n2285 VSS VSS nmos w=1u l=1u
M327 net91 n2286 VSS VSS nmos w=1u l=1u
M328 net91 n2286 net92 VDD pmos w=2u l=1u
M329 n2284 net91 VDD VDD pmos w=2u l=1u
M330 net92 n2285 VDD VDD pmos w=2u l=1u
M331 n2247 n2286 net93 VSS nmos w=1u l=1u
M332 net93 n2285 VSS VSS nmos w=1u l=1u
M333 n2247 n2286 VDD VDD pmos w=2u l=1u
M334 n2247 n2285 VDD VDD pmos w=2u l=1u
M335 n2286 n2288 net94 VSS nmos w=1u l=1u
M336 net94 n2287 VSS VSS nmos w=1u l=1u
M337 n2286 n2288 VDD VDD pmos w=2u l=1u
M338 n2286 n2287 VDD VDD pmos w=2u l=1u
M339 n2287 n2290 net95 VSS nmos w=1u l=1u
M340 net95 n2289 VSS VSS nmos w=1u l=1u
M341 n2287 n2290 VDD VDD pmos w=2u l=1u
M342 n2287 n2289 VDD VDD pmos w=2u l=1u
M343 net96 n2249 VSS VSS nmos w=1u l=1u
M344 net97 n2248 VSS VSS nmos w=1u l=1u
M345 n2285 net98 VSS VSS nmos w=1u l=1u
M346 net98 n2249 net99 VSS nmos w=1u l=1u
M347 net98 net96 net97 VSS nmos w=1u l=1u
M348 net99 net97 VSS VSS nmos w=1u l=1u
M349 net98 net96 net100 VDD pmos w=2u l=1u
M350 net96 n2249 VDD VDD pmos w=2u l=1u
M351 net97 n2249 net98 VDD pmos w=2u l=1u
M352 net97 n2248 VDD VDD pmos w=2u l=1u
M353 n2285 net98 VDD VDD pmos w=2u l=1u
M354 net100 net97 VDD VDD pmos w=2u l=1u
M355 n2249 n2292 net101 VSS nmos w=1u l=1u
M356 net101 n2291 VSS VSS nmos w=1u l=1u
M357 n2249 n2292 VDD VDD pmos w=2u l=1u
M358 n2249 n2291 VDD VDD pmos w=2u l=1u
M359 n2291 n2294 net102 VSS nmos w=1u l=1u
M360 net102 n2293 VSS VSS nmos w=1u l=1u
M361 n2291 n2294 VDD VDD pmos w=2u l=1u
M362 n2291 n2293 VDD VDD pmos w=2u l=1u
M363 net103 n2282 VSS VSS nmos w=1u l=1u
M364 net104 n2283 VSS VSS nmos w=1u l=1u
M365 n2248 net105 VSS VSS nmos w=1u l=1u
M366 net105 n2282 net106 VSS nmos w=1u l=1u
M367 net105 net103 net104 VSS nmos w=1u l=1u
M368 net106 net104 VSS VSS nmos w=1u l=1u
M369 net105 net103 net107 VDD pmos w=2u l=1u
M370 net103 n2282 VDD VDD pmos w=2u l=1u
M371 net104 n2282 net105 VDD pmos w=2u l=1u
M372 net104 n2283 VDD VDD pmos w=2u l=1u
M373 n2248 net105 VDD VDD pmos w=2u l=1u
M374 net107 net104 VDD VDD pmos w=2u l=1u
M375 n2282 net108 VSS VSS nmos w=1u l=1u
M376 net109 n2281 VSS VSS nmos w=1u l=1u
M377 net108 n2295 net109 VSS nmos w=1u l=1u
M378 net108 n2281 VDD VDD pmos w=2u l=1u
M379 net108 n2295 VDD VDD pmos w=2u l=1u
M380 n2282 net108 VDD VDD pmos w=2u l=1u
M381 n2281 n2297 net110 VSS nmos w=1u l=1u
M382 net110 n2296 VSS VSS nmos w=1u l=1u
M383 n2281 n2297 VDD VDD pmos w=2u l=1u
M384 n2281 n2296 VDD VDD pmos w=2u l=1u
M385 n2297 n2299 net111 VSS nmos w=1u l=1u
M386 net111 n2298 VSS VSS nmos w=1u l=1u
M387 n2297 n2299 VDD VDD pmos w=2u l=1u
M388 n2297 n2298 VDD VDD pmos w=2u l=1u
M389 n2298 net112 VSS VSS nmos w=1u l=1u
M390 net112 n2300 VSS VSS nmos w=1u l=1u
M391 net112 n2301 VSS VSS nmos w=1u l=1u
M392 net112 n2301 net113 VDD pmos w=2u l=1u
M393 n2298 net112 VDD VDD pmos w=2u l=1u
M394 net113 n2300 VDD VDD pmos w=2u l=1u
M395 net114 n2260 VSS VSS nmos w=1u l=1u
M396 net115 n2261 VSS VSS nmos w=1u l=1u
M397 n2296 net116 VSS VSS nmos w=1u l=1u
M398 net116 n2260 net117 VSS nmos w=1u l=1u
M399 net116 net114 net115 VSS nmos w=1u l=1u
M400 net117 net115 VSS VSS nmos w=1u l=1u
M401 net116 net114 net118 VDD pmos w=2u l=1u
M402 net114 n2260 VDD VDD pmos w=2u l=1u
M403 net115 n2260 net116 VDD pmos w=2u l=1u
M404 net115 n2261 VDD VDD pmos w=2u l=1u
M405 n2296 net116 VDD VDD pmos w=2u l=1u
M406 net118 net115 VDD VDD pmos w=2u l=1u
M407 n2260 n2302 VDD VDD pmos w=2u l=1u
M408 n2260 n2302 VSS VSS nmos w=1u l=1u
M409 n2295 n2304 net119 VSS nmos w=1u l=1u
M410 net119 n2303 VSS VSS nmos w=1u l=1u
M411 n2295 n2304 VDD VDD pmos w=2u l=1u
M412 n2295 n2303 VDD VDD pmos w=2u l=1u
M413 net120 n2261 VSS VSS nmos w=1u l=1u
M414 net121 n2302 VSS VSS nmos w=1u l=1u
M415 n2304 net122 VSS VSS nmos w=1u l=1u
M416 net122 n2261 net123 VSS nmos w=1u l=1u
M417 net122 net120 net121 VSS nmos w=1u l=1u
M418 net123 net121 VSS VSS nmos w=1u l=1u
M419 net122 net120 net124 VDD pmos w=2u l=1u
M420 net120 n2261 VDD VDD pmos w=2u l=1u
M421 net121 n2261 net122 VDD pmos w=2u l=1u
M422 net121 n2302 VDD VDD pmos w=2u l=1u
M423 n2304 net122 VDD VDD pmos w=2u l=1u
M424 net124 net121 VDD VDD pmos w=2u l=1u
M425 n2261 N511 net125 VSS nmos w=1u l=1u
M426 net125 N222 VSS VSS nmos w=1u l=1u
M427 n2261 N511 VDD VDD pmos w=2u l=1u
M428 n2261 N222 VDD VDD pmos w=2u l=1u
M429 n2302 n2258 net126 VSS nmos w=1u l=1u
M430 net126 n2305 VSS VSS nmos w=1u l=1u
M431 n2302 n2258 VDD VDD pmos w=2u l=1u
M432 n2302 n2305 VDD VDD pmos w=2u l=1u
M433 n2258 n2307 net127 VSS nmos w=1u l=1u
M434 net127 n2306 VSS VSS nmos w=1u l=1u
M435 n2258 n2307 VDD VDD pmos w=2u l=1u
M436 n2258 n2306 VDD VDD pmos w=2u l=1u
M437 n2307 n2309 net128 VSS nmos w=1u l=1u
M438 net128 n2308 VSS VSS nmos w=1u l=1u
M439 n2307 n2309 VDD VDD pmos w=2u l=1u
M440 n2307 n2308 VDD VDD pmos w=2u l=1u
M441 n2305 n2308 net129 VSS nmos w=1u l=1u
M442 net129 n2310 VSS VSS nmos w=1u l=1u
M443 n2305 n2308 VDD VDD pmos w=2u l=1u
M444 n2305 n2310 VDD VDD pmos w=2u l=1u
M445 n2308 n2312 net130 VSS nmos w=1u l=1u
M446 net130 n2311 VSS VSS nmos w=1u l=1u
M447 n2308 n2312 VDD VDD pmos w=2u l=1u
M448 n2308 n2311 VDD VDD pmos w=2u l=1u
M449 n2310 n2306 VSS VSS nmos w=1u l=1u
M450 n2310 n2313 VSS VSS nmos w=1u l=1u
M451 n2310 n2306 net131 VDD pmos w=2u l=1u
M452 net131 n2313 VDD VDD pmos w=2u l=1u
M453 n2306 net132 VSS VSS nmos w=1u l=1u
M454 net133 n2314 VSS VSS nmos w=1u l=1u
M455 net132 n2276 net133 VSS nmos w=1u l=1u
M456 net132 n2314 VDD VDD pmos w=2u l=1u
M457 net132 n2276 VDD VDD pmos w=2u l=1u
M458 n2306 net132 VDD VDD pmos w=2u l=1u
M459 n2314 N494 net134 VSS nmos w=1u l=1u
M460 net134 n2315 VSS VSS nmos w=1u l=1u
M461 n2314 N494 VDD VDD pmos w=2u l=1u
M462 n2314 n2315 VDD VDD pmos w=2u l=1u
M463 n2315 n2317 VSS VSS nmos w=1u l=1u
M464 n2315 n2316 VSS VSS nmos w=1u l=1u
M465 n2315 n2317 net135 VDD pmos w=2u l=1u
M466 net135 n2316 VDD VDD pmos w=2u l=1u
M467 n2317 n2319 VSS VSS nmos w=1u l=1u
M468 n2317 n2318 VSS VSS nmos w=1u l=1u
M469 n2317 n2319 net136 VDD pmos w=2u l=1u
M470 net136 n2318 VDD VDD pmos w=2u l=1u
M471 n2319 n2270 net137 VSS nmos w=1u l=1u
M472 net137 n2320 VSS VSS nmos w=1u l=1u
M473 n2319 n2270 VDD VDD pmos w=2u l=1u
M474 n2319 n2320 VDD VDD pmos w=2u l=1u
M475 n2320 n2321 net138 VSS nmos w=1u l=1u
M476 net138 N239 VSS VSS nmos w=1u l=1u
M477 n2320 n2321 VDD VDD pmos w=2u l=1u
M478 n2320 N239 VDD VDD pmos w=2u l=1u
M479 n2318 n2279 VDD VDD pmos w=2u l=1u
M480 n2318 n2279 VSS VSS nmos w=1u l=1u
M481 n2316 n2279 VSS VSS nmos w=1u l=1u
M482 n2316 N477 VSS VSS nmos w=1u l=1u
M483 n2316 n2279 net139 VDD pmos w=2u l=1u
M484 net139 N477 VDD VDD pmos w=2u l=1u
M485 n2276 n2323 net140 VSS nmos w=1u l=1u
M486 net140 n2322 VSS VSS nmos w=1u l=1u
M487 n2276 n2323 VDD VDD pmos w=2u l=1u
M488 n2276 n2322 VDD VDD pmos w=2u l=1u
M489 n2323 N239 net141 VSS nmos w=1u l=1u
M490 net141 N494 VSS VSS nmos w=1u l=1u
M491 n2323 N239 VDD VDD pmos w=2u l=1u
M492 n2323 N494 VDD VDD pmos w=2u l=1u
M493 net142 n2278 VSS VSS nmos w=1u l=1u
M494 net143 n2279 VSS VSS nmos w=1u l=1u
M495 n2322 net144 VSS VSS nmos w=1u l=1u
M496 net144 n2278 net145 VSS nmos w=1u l=1u
M497 net144 net142 net143 VSS nmos w=1u l=1u
M498 net145 net143 VSS VSS nmos w=1u l=1u
M499 net144 net142 net146 VDD pmos w=2u l=1u
M500 net142 n2278 VDD VDD pmos w=2u l=1u
M501 net143 n2278 net144 VDD pmos w=2u l=1u
M502 net143 n2279 VDD VDD pmos w=2u l=1u
M503 n2322 net144 VDD VDD pmos w=2u l=1u
M504 net146 net143 VDD VDD pmos w=2u l=1u
M505 n2278 N256 net147 VSS nmos w=1u l=1u
M506 net147 N477 VSS VSS nmos w=1u l=1u
M507 n2278 N256 VDD VDD pmos w=2u l=1u
M508 n2278 N477 VDD VDD pmos w=2u l=1u
M509 n2279 n2325 net148 VSS nmos w=1u l=1u
M510 net148 n2324 VSS VSS nmos w=1u l=1u
M511 n2279 n2325 VDD VDD pmos w=2u l=1u
M512 n2279 n2324 VDD VDD pmos w=2u l=1u
M513 n2325 n2327 net149 VSS nmos w=1u l=1u
M514 net149 n2326 VSS VSS nmos w=1u l=1u
M515 n2325 n2327 VDD VDD pmos w=2u l=1u
M516 n2325 n2326 VDD VDD pmos w=2u l=1u
M517 n2313 n2309 VDD VDD pmos w=2u l=1u
M518 n2313 n2309 VSS VSS nmos w=1u l=1u
M519 n2303 n2329 VSS VSS nmos w=1u l=1u
M520 n2303 n2328 VSS VSS nmos w=1u l=1u
M521 n2303 n2329 net150 VDD pmos w=2u l=1u
M522 net150 n2328 VDD VDD pmos w=2u l=1u
M523 n2329 n2300 VSS VSS nmos w=1u l=1u
M524 n2329 n2301 VSS VSS nmos w=1u l=1u
M525 n2329 n2300 net151 VDD pmos w=2u l=1u
M526 net151 n2301 VDD VDD pmos w=2u l=1u
M527 n2328 n2299 VDD VDD pmos w=2u l=1u
M528 n2328 n2299 VSS VSS nmos w=1u l=1u
M529 n2283 N528 net152 VSS nmos w=1u l=1u
M530 net152 N205 VSS VSS nmos w=1u l=1u
M531 n2283 N528 VDD VDD pmos w=2u l=1u
M532 n2283 N205 VDD VDD pmos w=2u l=1u
M533 N6250 n2330 net153 VSS nmos w=1u l=1u
M534 net153 n2288 VSS VSS nmos w=1u l=1u
M535 N6250 n2330 VDD VDD pmos w=2u l=1u
M536 N6250 n2288 VDD VDD pmos w=2u l=1u
M537 n2330 net154 VSS VSS nmos w=1u l=1u
M538 net154 n2331 VSS VSS nmos w=1u l=1u
M539 net154 n2332 VSS VSS nmos w=1u l=1u
M540 net154 n2332 net155 VDD pmos w=2u l=1u
M541 n2330 net154 VDD VDD pmos w=2u l=1u
M542 net155 n2331 VDD VDD pmos w=2u l=1u
M543 n2288 n2332 net156 VSS nmos w=1u l=1u
M544 net156 n2331 VSS VSS nmos w=1u l=1u
M545 n2288 n2332 VDD VDD pmos w=2u l=1u
M546 n2288 n2331 VDD VDD pmos w=2u l=1u
M547 n2332 n2334 net157 VSS nmos w=1u l=1u
M548 net157 n2333 VSS VSS nmos w=1u l=1u
M549 n2332 n2334 VDD VDD pmos w=2u l=1u
M550 n2332 n2333 VDD VDD pmos w=2u l=1u
M551 n2333 n2336 net158 VSS nmos w=1u l=1u
M552 net158 n2335 VSS VSS nmos w=1u l=1u
M553 n2333 n2336 VDD VDD pmos w=2u l=1u
M554 n2333 n2335 VDD VDD pmos w=2u l=1u
M555 net159 n2290 VSS VSS nmos w=1u l=1u
M556 net160 n2289 VSS VSS nmos w=1u l=1u
M557 n2331 net161 VSS VSS nmos w=1u l=1u
M558 net161 n2290 net162 VSS nmos w=1u l=1u
M559 net161 net159 net160 VSS nmos w=1u l=1u
M560 net162 net160 VSS VSS nmos w=1u l=1u
M561 net161 net159 net163 VDD pmos w=2u l=1u
M562 net159 n2290 VDD VDD pmos w=2u l=1u
M563 net160 n2290 net161 VDD pmos w=2u l=1u
M564 net160 n2289 VDD VDD pmos w=2u l=1u
M565 n2331 net161 VDD VDD pmos w=2u l=1u
M566 net163 net160 VDD VDD pmos w=2u l=1u
M567 n2290 n2338 net164 VSS nmos w=1u l=1u
M568 net164 n2337 VSS VSS nmos w=1u l=1u
M569 n2290 n2338 VDD VDD pmos w=2u l=1u
M570 n2290 n2337 VDD VDD pmos w=2u l=1u
M571 n2337 n2340 net165 VSS nmos w=1u l=1u
M572 net165 n2339 VSS VSS nmos w=1u l=1u
M573 n2337 n2340 VDD VDD pmos w=2u l=1u
M574 n2337 n2339 VDD VDD pmos w=2u l=1u
M575 net166 n2293 VSS VSS nmos w=1u l=1u
M576 net167 n2294 VSS VSS nmos w=1u l=1u
M577 n2289 net168 VSS VSS nmos w=1u l=1u
M578 net168 n2293 net169 VSS nmos w=1u l=1u
M579 net168 net166 net167 VSS nmos w=1u l=1u
M580 net169 net167 VSS VSS nmos w=1u l=1u
M581 net168 net166 net170 VDD pmos w=2u l=1u
M582 net166 n2293 VDD VDD pmos w=2u l=1u
M583 net167 n2293 net168 VDD pmos w=2u l=1u
M584 net167 n2294 VDD VDD pmos w=2u l=1u
M585 n2289 net168 VDD VDD pmos w=2u l=1u
M586 net170 net167 VDD VDD pmos w=2u l=1u
M587 n2293 net171 VSS VSS nmos w=1u l=1u
M588 net172 n2292 VSS VSS nmos w=1u l=1u
M589 net171 n2341 net172 VSS nmos w=1u l=1u
M590 net171 n2292 VDD VDD pmos w=2u l=1u
M591 net171 n2341 VDD VDD pmos w=2u l=1u
M592 n2293 net171 VDD VDD pmos w=2u l=1u
M593 n2292 n2343 net173 VSS nmos w=1u l=1u
M594 net173 n2342 VSS VSS nmos w=1u l=1u
M595 n2292 n2343 VDD VDD pmos w=2u l=1u
M596 n2292 n2342 VDD VDD pmos w=2u l=1u
M597 n2343 n2345 net174 VSS nmos w=1u l=1u
M598 net174 n2344 VSS VSS nmos w=1u l=1u
M599 n2343 n2345 VDD VDD pmos w=2u l=1u
M600 n2343 n2344 VDD VDD pmos w=2u l=1u
M601 n2344 net175 VSS VSS nmos w=1u l=1u
M602 net175 n2346 VSS VSS nmos w=1u l=1u
M603 net175 n2347 VSS VSS nmos w=1u l=1u
M604 net175 n2347 net176 VDD pmos w=2u l=1u
M605 n2344 net175 VDD VDD pmos w=2u l=1u
M606 net176 n2346 VDD VDD pmos w=2u l=1u
M607 net177 n2300 VSS VSS nmos w=1u l=1u
M608 net178 n2301 VSS VSS nmos w=1u l=1u
M609 n2342 net179 VSS VSS nmos w=1u l=1u
M610 net179 n2300 net180 VSS nmos w=1u l=1u
M611 net179 net177 net178 VSS nmos w=1u l=1u
M612 net180 net178 VSS VSS nmos w=1u l=1u
M613 net179 net177 net181 VDD pmos w=2u l=1u
M614 net177 n2300 VDD VDD pmos w=2u l=1u
M615 net178 n2300 net179 VDD pmos w=2u l=1u
M616 net178 n2301 VDD VDD pmos w=2u l=1u
M617 n2342 net179 VDD VDD pmos w=2u l=1u
M618 net181 net178 VDD VDD pmos w=2u l=1u
M619 n2301 n2348 VDD VDD pmos w=2u l=1u
M620 n2301 n2348 VSS VSS nmos w=1u l=1u
M621 n2341 n2350 net182 VSS nmos w=1u l=1u
M622 net182 n2349 VSS VSS nmos w=1u l=1u
M623 n2341 n2350 VDD VDD pmos w=2u l=1u
M624 n2341 n2349 VDD VDD pmos w=2u l=1u
M625 net183 n2348 VSS VSS nmos w=1u l=1u
M626 net184 n2300 VSS VSS nmos w=1u l=1u
M627 n2350 net185 VSS VSS nmos w=1u l=1u
M628 net185 n2348 net186 VSS nmos w=1u l=1u
M629 net185 net183 net184 VSS nmos w=1u l=1u
M630 net186 net184 VSS VSS nmos w=1u l=1u
M631 net185 net183 net187 VDD pmos w=2u l=1u
M632 net183 n2348 VDD VDD pmos w=2u l=1u
M633 net184 n2348 net185 VDD pmos w=2u l=1u
M634 net184 n2300 VDD VDD pmos w=2u l=1u
M635 n2350 net185 VDD VDD pmos w=2u l=1u
M636 net187 net184 VDD VDD pmos w=2u l=1u
M637 n2348 N511 net188 VSS nmos w=1u l=1u
M638 net188 N205 VSS VSS nmos w=1u l=1u
M639 n2348 N511 VDD VDD pmos w=2u l=1u
M640 n2348 N205 VDD VDD pmos w=2u l=1u
M641 n2300 n2299 net189 VSS nmos w=1u l=1u
M642 net189 n2351 VSS VSS nmos w=1u l=1u
M643 n2300 n2299 VDD VDD pmos w=2u l=1u
M644 n2300 n2351 VDD VDD pmos w=2u l=1u
M645 n2299 n2353 net190 VSS nmos w=1u l=1u
M646 net190 n2352 VSS VSS nmos w=1u l=1u
M647 n2299 n2353 VDD VDD pmos w=2u l=1u
M648 n2299 n2352 VDD VDD pmos w=2u l=1u
M649 n2353 n2355 net191 VSS nmos w=1u l=1u
M650 net191 n2354 VSS VSS nmos w=1u l=1u
M651 n2353 n2355 VDD VDD pmos w=2u l=1u
M652 n2353 n2354 VDD VDD pmos w=2u l=1u
M653 n2354 n2357 net192 VSS nmos w=1u l=1u
M654 net192 n2356 VSS VSS nmos w=1u l=1u
M655 n2354 n2357 VDD VDD pmos w=2u l=1u
M656 n2354 n2356 VDD VDD pmos w=2u l=1u
M657 net193 n2311 VSS VSS nmos w=1u l=1u
M658 net194 n2312 VSS VSS nmos w=1u l=1u
M659 n2352 net195 VSS VSS nmos w=1u l=1u
M660 net195 n2311 net196 VSS nmos w=1u l=1u
M661 net195 net193 net194 VSS nmos w=1u l=1u
M662 net196 net194 VSS VSS nmos w=1u l=1u
M663 net195 net193 net197 VDD pmos w=2u l=1u
M664 net193 n2311 VDD VDD pmos w=2u l=1u
M665 net194 n2311 net195 VDD pmos w=2u l=1u
M666 net194 n2312 VDD VDD pmos w=2u l=1u
M667 n2352 net195 VDD VDD pmos w=2u l=1u
M668 net197 net194 VDD VDD pmos w=2u l=1u
M669 n2311 n2358 VDD VDD pmos w=2u l=1u
M670 n2311 n2358 VSS VSS nmos w=1u l=1u
M671 n2351 n2360 net198 VSS nmos w=1u l=1u
M672 net198 n2359 VSS VSS nmos w=1u l=1u
M673 n2351 n2360 VDD VDD pmos w=2u l=1u
M674 n2351 n2359 VDD VDD pmos w=2u l=1u
M675 net199 n2312 VSS VSS nmos w=1u l=1u
M676 net200 n2358 VSS VSS nmos w=1u l=1u
M677 n2360 net201 VSS VSS nmos w=1u l=1u
M678 net201 n2312 net202 VSS nmos w=1u l=1u
M679 net201 net199 net200 VSS nmos w=1u l=1u
M680 net202 net200 VSS VSS nmos w=1u l=1u
M681 net201 net199 net203 VDD pmos w=2u l=1u
M682 net199 n2312 VDD VDD pmos w=2u l=1u
M683 net200 n2312 net201 VDD pmos w=2u l=1u
M684 net200 n2358 VDD VDD pmos w=2u l=1u
M685 n2360 net201 VDD VDD pmos w=2u l=1u
M686 net203 net200 VDD VDD pmos w=2u l=1u
M687 n2312 N494 net204 VSS nmos w=1u l=1u
M688 net204 N222 VSS VSS nmos w=1u l=1u
M689 n2312 N494 VDD VDD pmos w=2u l=1u
M690 n2312 N222 VDD VDD pmos w=2u l=1u
M691 n2358 n2309 net205 VSS nmos w=1u l=1u
M692 net205 n2361 VSS VSS nmos w=1u l=1u
M693 n2358 n2309 VDD VDD pmos w=2u l=1u
M694 n2358 n2361 VDD VDD pmos w=2u l=1u
M695 n2309 n2363 net206 VSS nmos w=1u l=1u
M696 net206 n2362 VSS VSS nmos w=1u l=1u
M697 n2309 n2363 VDD VDD pmos w=2u l=1u
M698 n2309 n2362 VDD VDD pmos w=2u l=1u
M699 n2363 n2365 net207 VSS nmos w=1u l=1u
M700 net207 n2364 VSS VSS nmos w=1u l=1u
M701 n2363 n2365 VDD VDD pmos w=2u l=1u
M702 n2363 n2364 VDD VDD pmos w=2u l=1u
M703 n2361 n2364 net208 VSS nmos w=1u l=1u
M704 net208 n2366 VSS VSS nmos w=1u l=1u
M705 n2361 n2364 VDD VDD pmos w=2u l=1u
M706 n2361 n2366 VDD VDD pmos w=2u l=1u
M707 n2364 n2368 net209 VSS nmos w=1u l=1u
M708 net209 n2367 VSS VSS nmos w=1u l=1u
M709 n2364 n2368 VDD VDD pmos w=2u l=1u
M710 n2364 n2367 VDD VDD pmos w=2u l=1u
M711 n2366 n2362 VSS VSS nmos w=1u l=1u
M712 n2366 n2369 VSS VSS nmos w=1u l=1u
M713 n2366 n2362 net210 VDD pmos w=2u l=1u
M714 net210 n2369 VDD VDD pmos w=2u l=1u
M715 n2362 net211 VSS VSS nmos w=1u l=1u
M716 net212 n2370 VSS VSS nmos w=1u l=1u
M717 net211 n2324 net212 VSS nmos w=1u l=1u
M718 net211 n2370 VDD VDD pmos w=2u l=1u
M719 net211 n2324 VDD VDD pmos w=2u l=1u
M720 n2362 net211 VDD VDD pmos w=2u l=1u
M721 n2370 N477 net213 VSS nmos w=1u l=1u
M722 net213 n2371 VSS VSS nmos w=1u l=1u
M723 n2370 N477 VDD VDD pmos w=2u l=1u
M724 n2370 n2371 VDD VDD pmos w=2u l=1u
M725 n2371 n2373 VSS VSS nmos w=1u l=1u
M726 n2371 n2372 VSS VSS nmos w=1u l=1u
M727 n2371 n2373 net214 VDD pmos w=2u l=1u
M728 net214 n2372 VDD VDD pmos w=2u l=1u
M729 n2373 n2375 VSS VSS nmos w=1u l=1u
M730 n2373 n2374 VSS VSS nmos w=1u l=1u
M731 n2373 n2375 net215 VDD pmos w=2u l=1u
M732 net215 n2374 VDD VDD pmos w=2u l=1u
M733 n2375 n2270 net216 VSS nmos w=1u l=1u
M734 net216 n2376 VSS VSS nmos w=1u l=1u
M735 n2375 n2270 VDD VDD pmos w=2u l=1u
M736 n2375 n2376 VDD VDD pmos w=2u l=1u
M737 n2376 n2377 net217 VSS nmos w=1u l=1u
M738 net217 N239 VSS VSS nmos w=1u l=1u
M739 n2376 n2377 VDD VDD pmos w=2u l=1u
M740 n2376 N239 VDD VDD pmos w=2u l=1u
M741 n2374 n2327 VDD VDD pmos w=2u l=1u
M742 n2374 n2327 VSS VSS nmos w=1u l=1u
M743 n2372 n2327 VSS VSS nmos w=1u l=1u
M744 n2372 N460 VSS VSS nmos w=1u l=1u
M745 n2372 n2327 net218 VDD pmos w=2u l=1u
M746 net218 N460 VDD VDD pmos w=2u l=1u
M747 n2324 n2379 net219 VSS nmos w=1u l=1u
M748 net219 n2378 VSS VSS nmos w=1u l=1u
M749 n2324 n2379 VDD VDD pmos w=2u l=1u
M750 n2324 n2378 VDD VDD pmos w=2u l=1u
M751 n2379 N239 net220 VSS nmos w=1u l=1u
M752 net220 N477 VSS VSS nmos w=1u l=1u
M753 n2379 N239 VDD VDD pmos w=2u l=1u
M754 n2379 N477 VDD VDD pmos w=2u l=1u
M755 net221 n2326 VSS VSS nmos w=1u l=1u
M756 net222 n2327 VSS VSS nmos w=1u l=1u
M757 n2378 net223 VSS VSS nmos w=1u l=1u
M758 net223 n2326 net224 VSS nmos w=1u l=1u
M759 net223 net221 net222 VSS nmos w=1u l=1u
M760 net224 net222 VSS VSS nmos w=1u l=1u
M761 net223 net221 net225 VDD pmos w=2u l=1u
M762 net221 n2326 VDD VDD pmos w=2u l=1u
M763 net222 n2326 net223 VDD pmos w=2u l=1u
M764 net222 n2327 VDD VDD pmos w=2u l=1u
M765 n2378 net223 VDD VDD pmos w=2u l=1u
M766 net225 net222 VDD VDD pmos w=2u l=1u
M767 n2326 N256 net226 VSS nmos w=1u l=1u
M768 net226 N460 VSS VSS nmos w=1u l=1u
M769 n2326 N256 VDD VDD pmos w=2u l=1u
M770 n2326 N460 VDD VDD pmos w=2u l=1u
M771 n2327 n2381 net227 VSS nmos w=1u l=1u
M772 net227 n2380 VSS VSS nmos w=1u l=1u
M773 n2327 n2381 VDD VDD pmos w=2u l=1u
M774 n2327 n2380 VDD VDD pmos w=2u l=1u
M775 n2381 n2383 net228 VSS nmos w=1u l=1u
M776 net228 n2382 VSS VSS nmos w=1u l=1u
M777 n2381 n2383 VDD VDD pmos w=2u l=1u
M778 n2381 n2382 VDD VDD pmos w=2u l=1u
M779 n2369 n2365 VDD VDD pmos w=2u l=1u
M780 n2369 n2365 VSS VSS nmos w=1u l=1u
M781 n2359 n2385 VSS VSS nmos w=1u l=1u
M782 n2359 n2384 VSS VSS nmos w=1u l=1u
M783 n2359 n2385 net229 VDD pmos w=2u l=1u
M784 net229 n2384 VDD VDD pmos w=2u l=1u
M785 n2385 net230 VSS VSS nmos w=1u l=1u
M786 net231 n2356 VSS VSS nmos w=1u l=1u
M787 net230 n2357 net231 VSS nmos w=1u l=1u
M788 net230 n2356 VDD VDD pmos w=2u l=1u
M789 net230 n2357 VDD VDD pmos w=2u l=1u
M790 n2385 net230 VDD VDD pmos w=2u l=1u
M791 n2384 n2355 VDD VDD pmos w=2u l=1u
M792 n2384 n2355 VSS VSS nmos w=1u l=1u
M793 n2349 n2387 VSS VSS nmos w=1u l=1u
M794 n2349 n2386 VSS VSS nmos w=1u l=1u
M795 n2349 n2387 net232 VDD pmos w=2u l=1u
M796 net232 n2386 VDD VDD pmos w=2u l=1u
M797 n2387 n2346 VSS VSS nmos w=1u l=1u
M798 n2387 n2347 VSS VSS nmos w=1u l=1u
M799 n2387 n2346 net233 VDD pmos w=2u l=1u
M800 net233 n2347 VDD VDD pmos w=2u l=1u
M801 n2386 n2345 VDD VDD pmos w=2u l=1u
M802 n2386 n2345 VSS VSS nmos w=1u l=1u
M803 n2294 N528 net234 VSS nmos w=1u l=1u
M804 net234 N188 VSS VSS nmos w=1u l=1u
M805 n2294 N528 VDD VDD pmos w=2u l=1u
M806 n2294 N188 VDD VDD pmos w=2u l=1u
M807 N6240 n2388 net235 VSS nmos w=1u l=1u
M808 net235 n2334 VSS VSS nmos w=1u l=1u
M809 N6240 n2388 VDD VDD pmos w=2u l=1u
M810 N6240 n2334 VDD VDD pmos w=2u l=1u
M811 n2388 net236 VSS VSS nmos w=1u l=1u
M812 net236 n2389 VSS VSS nmos w=1u l=1u
M813 net236 n2390 VSS VSS nmos w=1u l=1u
M814 net236 n2390 net237 VDD pmos w=2u l=1u
M815 n2388 net236 VDD VDD pmos w=2u l=1u
M816 net237 n2389 VDD VDD pmos w=2u l=1u
M817 n2334 n2390 net238 VSS nmos w=1u l=1u
M818 net238 n2389 VSS VSS nmos w=1u l=1u
M819 n2334 n2390 VDD VDD pmos w=2u l=1u
M820 n2334 n2389 VDD VDD pmos w=2u l=1u
M821 n2390 n2392 net239 VSS nmos w=1u l=1u
M822 net239 n2391 VSS VSS nmos w=1u l=1u
M823 n2390 n2392 VDD VDD pmos w=2u l=1u
M824 n2390 n2391 VDD VDD pmos w=2u l=1u
M825 n2391 n2394 net240 VSS nmos w=1u l=1u
M826 net240 n2393 VSS VSS nmos w=1u l=1u
M827 n2391 n2394 VDD VDD pmos w=2u l=1u
M828 n2391 n2393 VDD VDD pmos w=2u l=1u
M829 net241 n2336 VSS VSS nmos w=1u l=1u
M830 net242 n2335 VSS VSS nmos w=1u l=1u
M831 n2389 net243 VSS VSS nmos w=1u l=1u
M832 net243 n2336 net244 VSS nmos w=1u l=1u
M833 net243 net241 net242 VSS nmos w=1u l=1u
M834 net244 net242 VSS VSS nmos w=1u l=1u
M835 net243 net241 net245 VDD pmos w=2u l=1u
M836 net241 n2336 VDD VDD pmos w=2u l=1u
M837 net242 n2336 net243 VDD pmos w=2u l=1u
M838 net242 n2335 VDD VDD pmos w=2u l=1u
M839 n2389 net243 VDD VDD pmos w=2u l=1u
M840 net245 net242 VDD VDD pmos w=2u l=1u
M841 n2336 n2396 net246 VSS nmos w=1u l=1u
M842 net246 n2395 VSS VSS nmos w=1u l=1u
M843 n2336 n2396 VDD VDD pmos w=2u l=1u
M844 n2336 n2395 VDD VDD pmos w=2u l=1u
M845 n2395 n2398 net247 VSS nmos w=1u l=1u
M846 net247 n2397 VSS VSS nmos w=1u l=1u
M847 n2395 n2398 VDD VDD pmos w=2u l=1u
M848 n2395 n2397 VDD VDD pmos w=2u l=1u
M849 net248 n2339 VSS VSS nmos w=1u l=1u
M850 net249 n2340 VSS VSS nmos w=1u l=1u
M851 n2335 net250 VSS VSS nmos w=1u l=1u
M852 net250 n2339 net251 VSS nmos w=1u l=1u
M853 net250 net248 net249 VSS nmos w=1u l=1u
M854 net251 net249 VSS VSS nmos w=1u l=1u
M855 net250 net248 net252 VDD pmos w=2u l=1u
M856 net248 n2339 VDD VDD pmos w=2u l=1u
M857 net249 n2339 net250 VDD pmos w=2u l=1u
M858 net249 n2340 VDD VDD pmos w=2u l=1u
M859 n2335 net250 VDD VDD pmos w=2u l=1u
M860 net252 net249 VDD VDD pmos w=2u l=1u
M861 n2339 net253 VSS VSS nmos w=1u l=1u
M862 net254 n2338 VSS VSS nmos w=1u l=1u
M863 net253 n2399 net254 VSS nmos w=1u l=1u
M864 net253 n2338 VDD VDD pmos w=2u l=1u
M865 net253 n2399 VDD VDD pmos w=2u l=1u
M866 n2339 net253 VDD VDD pmos w=2u l=1u
M867 n2338 n2401 net255 VSS nmos w=1u l=1u
M868 net255 n2400 VSS VSS nmos w=1u l=1u
M869 n2338 n2401 VDD VDD pmos w=2u l=1u
M870 n2338 n2400 VDD VDD pmos w=2u l=1u
M871 n2401 n2403 net256 VSS nmos w=1u l=1u
M872 net256 n2402 VSS VSS nmos w=1u l=1u
M873 n2401 n2403 VDD VDD pmos w=2u l=1u
M874 n2401 n2402 VDD VDD pmos w=2u l=1u
M875 n2402 net257 VSS VSS nmos w=1u l=1u
M876 net257 n2404 VSS VSS nmos w=1u l=1u
M877 net257 n2405 VSS VSS nmos w=1u l=1u
M878 net257 n2405 net258 VDD pmos w=2u l=1u
M879 n2402 net257 VDD VDD pmos w=2u l=1u
M880 net258 n2404 VDD VDD pmos w=2u l=1u
M881 net259 n2346 VSS VSS nmos w=1u l=1u
M882 net260 n2347 VSS VSS nmos w=1u l=1u
M883 n2400 net261 VSS VSS nmos w=1u l=1u
M884 net261 n2346 net262 VSS nmos w=1u l=1u
M885 net261 net259 net260 VSS nmos w=1u l=1u
M886 net262 net260 VSS VSS nmos w=1u l=1u
M887 net261 net259 net263 VDD pmos w=2u l=1u
M888 net259 n2346 VDD VDD pmos w=2u l=1u
M889 net260 n2346 net261 VDD pmos w=2u l=1u
M890 net260 n2347 VDD VDD pmos w=2u l=1u
M891 n2400 net261 VDD VDD pmos w=2u l=1u
M892 net263 net260 VDD VDD pmos w=2u l=1u
M893 n2347 n2406 VDD VDD pmos w=2u l=1u
M894 n2347 n2406 VSS VSS nmos w=1u l=1u
M895 n2399 n2408 net264 VSS nmos w=1u l=1u
M896 net264 n2407 VSS VSS nmos w=1u l=1u
M897 n2399 n2408 VDD VDD pmos w=2u l=1u
M898 n2399 n2407 VDD VDD pmos w=2u l=1u
M899 net265 n2406 VSS VSS nmos w=1u l=1u
M900 net266 n2346 VSS VSS nmos w=1u l=1u
M901 n2408 net267 VSS VSS nmos w=1u l=1u
M902 net267 n2406 net268 VSS nmos w=1u l=1u
M903 net267 net265 net266 VSS nmos w=1u l=1u
M904 net268 net266 VSS VSS nmos w=1u l=1u
M905 net267 net265 net269 VDD pmos w=2u l=1u
M906 net265 n2406 VDD VDD pmos w=2u l=1u
M907 net266 n2406 net267 VDD pmos w=2u l=1u
M908 net266 n2346 VDD VDD pmos w=2u l=1u
M909 n2408 net267 VDD VDD pmos w=2u l=1u
M910 net269 net266 VDD VDD pmos w=2u l=1u
M911 n2406 N511 net270 VSS nmos w=1u l=1u
M912 net270 N188 VSS VSS nmos w=1u l=1u
M913 n2406 N511 VDD VDD pmos w=2u l=1u
M914 n2406 N188 VDD VDD pmos w=2u l=1u
M915 n2346 n2345 net271 VSS nmos w=1u l=1u
M916 net271 n2409 VSS VSS nmos w=1u l=1u
M917 n2346 n2345 VDD VDD pmos w=2u l=1u
M918 n2346 n2409 VDD VDD pmos w=2u l=1u
M919 n2345 n2411 net272 VSS nmos w=1u l=1u
M920 net272 n2410 VSS VSS nmos w=1u l=1u
M921 n2345 n2411 VDD VDD pmos w=2u l=1u
M922 n2345 n2410 VDD VDD pmos w=2u l=1u
M923 n2411 n2413 net273 VSS nmos w=1u l=1u
M924 net273 n2412 VSS VSS nmos w=1u l=1u
M925 n2411 n2413 VDD VDD pmos w=2u l=1u
M926 n2411 n2412 VDD VDD pmos w=2u l=1u
M927 n2412 net274 VSS VSS nmos w=1u l=1u
M928 net274 n2414 VSS VSS nmos w=1u l=1u
M929 net274 n2415 VSS VSS nmos w=1u l=1u
M930 net274 n2415 net275 VDD pmos w=2u l=1u
M931 n2412 net274 VDD VDD pmos w=2u l=1u
M932 net275 n2414 VDD VDD pmos w=2u l=1u
M933 net276 n2356 VSS VSS nmos w=1u l=1u
M934 net277 n2357 VSS VSS nmos w=1u l=1u
M935 n2410 net278 VSS VSS nmos w=1u l=1u
M936 net278 n2356 net279 VSS nmos w=1u l=1u
M937 net278 net276 net277 VSS nmos w=1u l=1u
M938 net279 net277 VSS VSS nmos w=1u l=1u
M939 net278 net276 net280 VDD pmos w=2u l=1u
M940 net276 n2356 VDD VDD pmos w=2u l=1u
M941 net277 n2356 net278 VDD pmos w=2u l=1u
M942 net277 n2357 VDD VDD pmos w=2u l=1u
M943 n2410 net278 VDD VDD pmos w=2u l=1u
M944 net280 net277 VDD VDD pmos w=2u l=1u
M945 n2356 n2416 VDD VDD pmos w=2u l=1u
M946 n2356 n2416 VSS VSS nmos w=1u l=1u
M947 n2409 n2418 net281 VSS nmos w=1u l=1u
M948 net281 n2417 VSS VSS nmos w=1u l=1u
M949 n2409 n2418 VDD VDD pmos w=2u l=1u
M950 n2409 n2417 VDD VDD pmos w=2u l=1u
M951 net282 n2357 VSS VSS nmos w=1u l=1u
M952 net283 n2416 VSS VSS nmos w=1u l=1u
M953 n2418 net284 VSS VSS nmos w=1u l=1u
M954 net284 n2357 net285 VSS nmos w=1u l=1u
M955 net284 net282 net283 VSS nmos w=1u l=1u
M956 net285 net283 VSS VSS nmos w=1u l=1u
M957 net284 net282 net286 VDD pmos w=2u l=1u
M958 net282 n2357 VDD VDD pmos w=2u l=1u
M959 net283 n2357 net284 VDD pmos w=2u l=1u
M960 net283 n2416 VDD VDD pmos w=2u l=1u
M961 n2418 net284 VDD VDD pmos w=2u l=1u
M962 net286 net283 VDD VDD pmos w=2u l=1u
M963 n2357 N494 net287 VSS nmos w=1u l=1u
M964 net287 N205 VSS VSS nmos w=1u l=1u
M965 n2357 N494 VDD VDD pmos w=2u l=1u
M966 n2357 N205 VDD VDD pmos w=2u l=1u
M967 n2416 n2355 net288 VSS nmos w=1u l=1u
M968 net288 n2419 VSS VSS nmos w=1u l=1u
M969 n2416 n2355 VDD VDD pmos w=2u l=1u
M970 n2416 n2419 VDD VDD pmos w=2u l=1u
M971 n2355 n2421 net289 VSS nmos w=1u l=1u
M972 net289 n2420 VSS VSS nmos w=1u l=1u
M973 n2355 n2421 VDD VDD pmos w=2u l=1u
M974 n2355 n2420 VDD VDD pmos w=2u l=1u
M975 n2421 n2423 net290 VSS nmos w=1u l=1u
M976 net290 n2422 VSS VSS nmos w=1u l=1u
M977 n2421 n2423 VDD VDD pmos w=2u l=1u
M978 n2421 n2422 VDD VDD pmos w=2u l=1u
M979 n2422 net291 VSS VSS nmos w=1u l=1u
M980 net291 n2424 VSS VSS nmos w=1u l=1u
M981 net291 n2425 VSS VSS nmos w=1u l=1u
M982 net291 n2425 net292 VDD pmos w=2u l=1u
M983 n2422 net291 VDD VDD pmos w=2u l=1u
M984 net292 n2424 VDD VDD pmos w=2u l=1u
M985 net293 n2367 VSS VSS nmos w=1u l=1u
M986 net294 n2368 VSS VSS nmos w=1u l=1u
M987 n2420 net295 VSS VSS nmos w=1u l=1u
M988 net295 n2367 net296 VSS nmos w=1u l=1u
M989 net295 net293 net294 VSS nmos w=1u l=1u
M990 net296 net294 VSS VSS nmos w=1u l=1u
M991 net295 net293 net297 VDD pmos w=2u l=1u
M992 net293 n2367 VDD VDD pmos w=2u l=1u
M993 net294 n2367 net295 VDD pmos w=2u l=1u
M994 net294 n2368 VDD VDD pmos w=2u l=1u
M995 n2420 net295 VDD VDD pmos w=2u l=1u
M996 net297 net294 VDD VDD pmos w=2u l=1u
M997 n2367 n2426 VDD VDD pmos w=2u l=1u
M998 n2367 n2426 VSS VSS nmos w=1u l=1u
M999 n2419 n2428 net298 VSS nmos w=1u l=1u
M1000 net298 n2427 VSS VSS nmos w=1u l=1u
M1001 n2419 n2428 VDD VDD pmos w=2u l=1u
M1002 n2419 n2427 VDD VDD pmos w=2u l=1u
M1003 net299 n2368 VSS VSS nmos w=1u l=1u
M1004 net300 n2426 VSS VSS nmos w=1u l=1u
M1005 n2428 net301 VSS VSS nmos w=1u l=1u
M1006 net301 n2368 net302 VSS nmos w=1u l=1u
M1007 net301 net299 net300 VSS nmos w=1u l=1u
M1008 net302 net300 VSS VSS nmos w=1u l=1u
M1009 net301 net299 net303 VDD pmos w=2u l=1u
M1010 net299 n2368 VDD VDD pmos w=2u l=1u
M1011 net300 n2368 net301 VDD pmos w=2u l=1u
M1012 net300 n2426 VDD VDD pmos w=2u l=1u
M1013 n2428 net301 VDD VDD pmos w=2u l=1u
M1014 net303 net300 VDD VDD pmos w=2u l=1u
M1015 n2368 N477 net304 VSS nmos w=1u l=1u
M1016 net304 N222 VSS VSS nmos w=1u l=1u
M1017 n2368 N477 VDD VDD pmos w=2u l=1u
M1018 n2368 N222 VDD VDD pmos w=2u l=1u
M1019 n2426 n2365 net305 VSS nmos w=1u l=1u
M1020 net305 n2429 VSS VSS nmos w=1u l=1u
M1021 n2426 n2365 VDD VDD pmos w=2u l=1u
M1022 n2426 n2429 VDD VDD pmos w=2u l=1u
M1023 n2365 n2431 net306 VSS nmos w=1u l=1u
M1024 net306 n2430 VSS VSS nmos w=1u l=1u
M1025 n2365 n2431 VDD VDD pmos w=2u l=1u
M1026 n2365 n2430 VDD VDD pmos w=2u l=1u
M1027 n2431 n2433 net307 VSS nmos w=1u l=1u
M1028 net307 n2432 VSS VSS nmos w=1u l=1u
M1029 n2431 n2433 VDD VDD pmos w=2u l=1u
M1030 n2431 n2432 VDD VDD pmos w=2u l=1u
M1031 n2429 n2432 net308 VSS nmos w=1u l=1u
M1032 net308 n2434 VSS VSS nmos w=1u l=1u
M1033 n2429 n2432 VDD VDD pmos w=2u l=1u
M1034 n2429 n2434 VDD VDD pmos w=2u l=1u
M1035 n2432 n2436 net309 VSS nmos w=1u l=1u
M1036 net309 n2435 VSS VSS nmos w=1u l=1u
M1037 n2432 n2436 VDD VDD pmos w=2u l=1u
M1038 n2432 n2435 VDD VDD pmos w=2u l=1u
M1039 n2434 n2430 VSS VSS nmos w=1u l=1u
M1040 n2434 n2437 VSS VSS nmos w=1u l=1u
M1041 n2434 n2430 net310 VDD pmos w=2u l=1u
M1042 net310 n2437 VDD VDD pmos w=2u l=1u
M1043 n2430 net311 VSS VSS nmos w=1u l=1u
M1044 net312 n2438 VSS VSS nmos w=1u l=1u
M1045 net311 n2380 net312 VSS nmos w=1u l=1u
M1046 net311 n2438 VDD VDD pmos w=2u l=1u
M1047 net311 n2380 VDD VDD pmos w=2u l=1u
M1048 n2430 net311 VDD VDD pmos w=2u l=1u
M1049 n2438 N460 net313 VSS nmos w=1u l=1u
M1050 net313 n2439 VSS VSS nmos w=1u l=1u
M1051 n2438 N460 VDD VDD pmos w=2u l=1u
M1052 n2438 n2439 VDD VDD pmos w=2u l=1u
M1053 n2439 n2441 VSS VSS nmos w=1u l=1u
M1054 n2439 n2440 VSS VSS nmos w=1u l=1u
M1055 n2439 n2441 net314 VDD pmos w=2u l=1u
M1056 net314 n2440 VDD VDD pmos w=2u l=1u
M1057 n2441 n2443 VSS VSS nmos w=1u l=1u
M1058 n2441 n2442 VSS VSS nmos w=1u l=1u
M1059 n2441 n2443 net315 VDD pmos w=2u l=1u
M1060 net315 n2442 VDD VDD pmos w=2u l=1u
M1061 n2443 n2270 net316 VSS nmos w=1u l=1u
M1062 net316 n2444 VSS VSS nmos w=1u l=1u
M1063 n2443 n2270 VDD VDD pmos w=2u l=1u
M1064 n2443 n2444 VDD VDD pmos w=2u l=1u
M1065 n2444 n2445 net317 VSS nmos w=1u l=1u
M1066 net317 N239 VSS VSS nmos w=1u l=1u
M1067 n2444 n2445 VDD VDD pmos w=2u l=1u
M1068 n2444 N239 VDD VDD pmos w=2u l=1u
M1069 n2442 n2383 VDD VDD pmos w=2u l=1u
M1070 n2442 n2383 VSS VSS nmos w=1u l=1u
M1071 n2440 n2383 VSS VSS nmos w=1u l=1u
M1072 n2440 N443 VSS VSS nmos w=1u l=1u
M1073 n2440 n2383 net318 VDD pmos w=2u l=1u
M1074 net318 N443 VDD VDD pmos w=2u l=1u
M1075 n2380 n2447 net319 VSS nmos w=1u l=1u
M1076 net319 n2446 VSS VSS nmos w=1u l=1u
M1077 n2380 n2447 VDD VDD pmos w=2u l=1u
M1078 n2380 n2446 VDD VDD pmos w=2u l=1u
M1079 n2447 N239 net320 VSS nmos w=1u l=1u
M1080 net320 N460 VSS VSS nmos w=1u l=1u
M1081 n2447 N239 VDD VDD pmos w=2u l=1u
M1082 n2447 N460 VDD VDD pmos w=2u l=1u
M1083 net321 n2382 VSS VSS nmos w=1u l=1u
M1084 net322 n2383 VSS VSS nmos w=1u l=1u
M1085 n2446 net323 VSS VSS nmos w=1u l=1u
M1086 net323 n2382 net324 VSS nmos w=1u l=1u
M1087 net323 net321 net322 VSS nmos w=1u l=1u
M1088 net324 net322 VSS VSS nmos w=1u l=1u
M1089 net323 net321 net325 VDD pmos w=2u l=1u
M1090 net321 n2382 VDD VDD pmos w=2u l=1u
M1091 net322 n2382 net323 VDD pmos w=2u l=1u
M1092 net322 n2383 VDD VDD pmos w=2u l=1u
M1093 n2446 net323 VDD VDD pmos w=2u l=1u
M1094 net325 net322 VDD VDD pmos w=2u l=1u
M1095 n2382 N256 net326 VSS nmos w=1u l=1u
M1096 net326 N443 VSS VSS nmos w=1u l=1u
M1097 n2382 N256 VDD VDD pmos w=2u l=1u
M1098 n2382 N443 VDD VDD pmos w=2u l=1u
M1099 n2383 n2449 net327 VSS nmos w=1u l=1u
M1100 net327 n2448 VSS VSS nmos w=1u l=1u
M1101 n2383 n2449 VDD VDD pmos w=2u l=1u
M1102 n2383 n2448 VDD VDD pmos w=2u l=1u
M1103 n2449 n2451 net328 VSS nmos w=1u l=1u
M1104 net328 n2450 VSS VSS nmos w=1u l=1u
M1105 n2449 n2451 VDD VDD pmos w=2u l=1u
M1106 n2449 n2450 VDD VDD pmos w=2u l=1u
M1107 n2437 n2433 VDD VDD pmos w=2u l=1u
M1108 n2437 n2433 VSS VSS nmos w=1u l=1u
M1109 n2427 n2453 VSS VSS nmos w=1u l=1u
M1110 n2427 n2452 VSS VSS nmos w=1u l=1u
M1111 n2427 n2453 net329 VDD pmos w=2u l=1u
M1112 net329 n2452 VDD VDD pmos w=2u l=1u
M1113 n2453 n2424 VSS VSS nmos w=1u l=1u
M1114 n2453 n2425 VSS VSS nmos w=1u l=1u
M1115 n2453 n2424 net330 VDD pmos w=2u l=1u
M1116 net330 n2425 VDD VDD pmos w=2u l=1u
M1117 n2452 n2423 VDD VDD pmos w=2u l=1u
M1118 n2452 n2423 VSS VSS nmos w=1u l=1u
M1119 n2417 n2455 VSS VSS nmos w=1u l=1u
M1120 n2417 n2454 VSS VSS nmos w=1u l=1u
M1121 n2417 n2455 net331 VDD pmos w=2u l=1u
M1122 net331 n2454 VDD VDD pmos w=2u l=1u
M1123 n2455 n2414 VSS VSS nmos w=1u l=1u
M1124 n2455 n2415 VSS VSS nmos w=1u l=1u
M1125 n2455 n2414 net332 VDD pmos w=2u l=1u
M1126 net332 n2415 VDD VDD pmos w=2u l=1u
M1127 n2454 n2413 VDD VDD pmos w=2u l=1u
M1128 n2454 n2413 VSS VSS nmos w=1u l=1u
M1129 n2407 n2457 VSS VSS nmos w=1u l=1u
M1130 n2407 n2456 VSS VSS nmos w=1u l=1u
M1131 n2407 n2457 net333 VDD pmos w=2u l=1u
M1132 net333 n2456 VDD VDD pmos w=2u l=1u
M1133 n2457 n2404 VSS VSS nmos w=1u l=1u
M1134 n2457 n2405 VSS VSS nmos w=1u l=1u
M1135 n2457 n2404 net334 VDD pmos w=2u l=1u
M1136 net334 n2405 VDD VDD pmos w=2u l=1u
M1137 n2456 n2403 VDD VDD pmos w=2u l=1u
M1138 n2456 n2403 VSS VSS nmos w=1u l=1u
M1139 n2340 N528 net335 VSS nmos w=1u l=1u
M1140 net335 N171 VSS VSS nmos w=1u l=1u
M1141 n2340 N528 VDD VDD pmos w=2u l=1u
M1142 n2340 N171 VDD VDD pmos w=2u l=1u
M1143 N6230 n2458 net336 VSS nmos w=1u l=1u
M1144 net336 n2392 VSS VSS nmos w=1u l=1u
M1145 N6230 n2458 VDD VDD pmos w=2u l=1u
M1146 N6230 n2392 VDD VDD pmos w=2u l=1u
M1147 n2458 net337 VSS VSS nmos w=1u l=1u
M1148 net337 n2459 VSS VSS nmos w=1u l=1u
M1149 net337 n2460 VSS VSS nmos w=1u l=1u
M1150 net337 n2460 net338 VDD pmos w=2u l=1u
M1151 n2458 net337 VDD VDD pmos w=2u l=1u
M1152 net338 n2459 VDD VDD pmos w=2u l=1u
M1153 n2392 n2460 net339 VSS nmos w=1u l=1u
M1154 net339 n2459 VSS VSS nmos w=1u l=1u
M1155 n2392 n2460 VDD VDD pmos w=2u l=1u
M1156 n2392 n2459 VDD VDD pmos w=2u l=1u
M1157 n2460 n2462 net340 VSS nmos w=1u l=1u
M1158 net340 n2461 VSS VSS nmos w=1u l=1u
M1159 n2460 n2462 VDD VDD pmos w=2u l=1u
M1160 n2460 n2461 VDD VDD pmos w=2u l=1u
M1161 n2461 n2464 net341 VSS nmos w=1u l=1u
M1162 net341 n2463 VSS VSS nmos w=1u l=1u
M1163 n2461 n2464 VDD VDD pmos w=2u l=1u
M1164 n2461 n2463 VDD VDD pmos w=2u l=1u
M1165 net342 n2394 VSS VSS nmos w=1u l=1u
M1166 net343 n2393 VSS VSS nmos w=1u l=1u
M1167 n2459 net344 VSS VSS nmos w=1u l=1u
M1168 net344 n2394 net345 VSS nmos w=1u l=1u
M1169 net344 net342 net343 VSS nmos w=1u l=1u
M1170 net345 net343 VSS VSS nmos w=1u l=1u
M1171 net344 net342 net346 VDD pmos w=2u l=1u
M1172 net342 n2394 VDD VDD pmos w=2u l=1u
M1173 net343 n2394 net344 VDD pmos w=2u l=1u
M1174 net343 n2393 VDD VDD pmos w=2u l=1u
M1175 n2459 net344 VDD VDD pmos w=2u l=1u
M1176 net346 net343 VDD VDD pmos w=2u l=1u
M1177 n2394 n2466 net347 VSS nmos w=1u l=1u
M1178 net347 n2465 VSS VSS nmos w=1u l=1u
M1179 n2394 n2466 VDD VDD pmos w=2u l=1u
M1180 n2394 n2465 VDD VDD pmos w=2u l=1u
M1181 n2465 n2468 net348 VSS nmos w=1u l=1u
M1182 net348 n2467 VSS VSS nmos w=1u l=1u
M1183 n2465 n2468 VDD VDD pmos w=2u l=1u
M1184 n2465 n2467 VDD VDD pmos w=2u l=1u
M1185 net349 n2397 VSS VSS nmos w=1u l=1u
M1186 net350 n2398 VSS VSS nmos w=1u l=1u
M1187 n2393 net351 VSS VSS nmos w=1u l=1u
M1188 net351 n2397 net352 VSS nmos w=1u l=1u
M1189 net351 net349 net350 VSS nmos w=1u l=1u
M1190 net352 net350 VSS VSS nmos w=1u l=1u
M1191 net351 net349 net353 VDD pmos w=2u l=1u
M1192 net349 n2397 VDD VDD pmos w=2u l=1u
M1193 net350 n2397 net351 VDD pmos w=2u l=1u
M1194 net350 n2398 VDD VDD pmos w=2u l=1u
M1195 n2393 net351 VDD VDD pmos w=2u l=1u
M1196 net353 net350 VDD VDD pmos w=2u l=1u
M1197 n2397 net354 VSS VSS nmos w=1u l=1u
M1198 net355 n2396 VSS VSS nmos w=1u l=1u
M1199 net354 n2469 net355 VSS nmos w=1u l=1u
M1200 net354 n2396 VDD VDD pmos w=2u l=1u
M1201 net354 n2469 VDD VDD pmos w=2u l=1u
M1202 n2397 net354 VDD VDD pmos w=2u l=1u
M1203 n2396 n2471 net356 VSS nmos w=1u l=1u
M1204 net356 n2470 VSS VSS nmos w=1u l=1u
M1205 n2396 n2471 VDD VDD pmos w=2u l=1u
M1206 n2396 n2470 VDD VDD pmos w=2u l=1u
M1207 n2471 n2473 net357 VSS nmos w=1u l=1u
M1208 net357 n2472 VSS VSS nmos w=1u l=1u
M1209 n2471 n2473 VDD VDD pmos w=2u l=1u
M1210 n2471 n2472 VDD VDD pmos w=2u l=1u
M1211 n2472 net358 VSS VSS nmos w=1u l=1u
M1212 net358 n2474 VSS VSS nmos w=1u l=1u
M1213 net358 n2475 VSS VSS nmos w=1u l=1u
M1214 net358 n2475 net359 VDD pmos w=2u l=1u
M1215 n2472 net358 VDD VDD pmos w=2u l=1u
M1216 net359 n2474 VDD VDD pmos w=2u l=1u
M1217 net360 n2404 VSS VSS nmos w=1u l=1u
M1218 net361 n2405 VSS VSS nmos w=1u l=1u
M1219 n2470 net362 VSS VSS nmos w=1u l=1u
M1220 net362 n2404 net363 VSS nmos w=1u l=1u
M1221 net362 net360 net361 VSS nmos w=1u l=1u
M1222 net363 net361 VSS VSS nmos w=1u l=1u
M1223 net362 net360 net364 VDD pmos w=2u l=1u
M1224 net360 n2404 VDD VDD pmos w=2u l=1u
M1225 net361 n2404 net362 VDD pmos w=2u l=1u
M1226 net361 n2405 VDD VDD pmos w=2u l=1u
M1227 n2470 net362 VDD VDD pmos w=2u l=1u
M1228 net364 net361 VDD VDD pmos w=2u l=1u
M1229 n2405 n2476 VDD VDD pmos w=2u l=1u
M1230 n2405 n2476 VSS VSS nmos w=1u l=1u
M1231 n2469 n2478 net365 VSS nmos w=1u l=1u
M1232 net365 n2477 VSS VSS nmos w=1u l=1u
M1233 n2469 n2478 VDD VDD pmos w=2u l=1u
M1234 n2469 n2477 VDD VDD pmos w=2u l=1u
M1235 net366 n2476 VSS VSS nmos w=1u l=1u
M1236 net367 n2404 VSS VSS nmos w=1u l=1u
M1237 n2478 net368 VSS VSS nmos w=1u l=1u
M1238 net368 n2476 net369 VSS nmos w=1u l=1u
M1239 net368 net366 net367 VSS nmos w=1u l=1u
M1240 net369 net367 VSS VSS nmos w=1u l=1u
M1241 net368 net366 net370 VDD pmos w=2u l=1u
M1242 net366 n2476 VDD VDD pmos w=2u l=1u
M1243 net367 n2476 net368 VDD pmos w=2u l=1u
M1244 net367 n2404 VDD VDD pmos w=2u l=1u
M1245 n2478 net368 VDD VDD pmos w=2u l=1u
M1246 net370 net367 VDD VDD pmos w=2u l=1u
M1247 n2476 N511 net371 VSS nmos w=1u l=1u
M1248 net371 N171 VSS VSS nmos w=1u l=1u
M1249 n2476 N511 VDD VDD pmos w=2u l=1u
M1250 n2476 N171 VDD VDD pmos w=2u l=1u
M1251 n2404 n2403 net372 VSS nmos w=1u l=1u
M1252 net372 n2479 VSS VSS nmos w=1u l=1u
M1253 n2404 n2403 VDD VDD pmos w=2u l=1u
M1254 n2404 n2479 VDD VDD pmos w=2u l=1u
M1255 n2403 n2481 net373 VSS nmos w=1u l=1u
M1256 net373 n2480 VSS VSS nmos w=1u l=1u
M1257 n2403 n2481 VDD VDD pmos w=2u l=1u
M1258 n2403 n2480 VDD VDD pmos w=2u l=1u
M1259 n2481 n2483 net374 VSS nmos w=1u l=1u
M1260 net374 n2482 VSS VSS nmos w=1u l=1u
M1261 n2481 n2483 VDD VDD pmos w=2u l=1u
M1262 n2481 n2482 VDD VDD pmos w=2u l=1u
M1263 n2482 net375 VSS VSS nmos w=1u l=1u
M1264 net375 n2484 VSS VSS nmos w=1u l=1u
M1265 net375 n2485 VSS VSS nmos w=1u l=1u
M1266 net375 n2485 net376 VDD pmos w=2u l=1u
M1267 n2482 net375 VDD VDD pmos w=2u l=1u
M1268 net376 n2484 VDD VDD pmos w=2u l=1u
M1269 net377 n2414 VSS VSS nmos w=1u l=1u
M1270 net378 n2415 VSS VSS nmos w=1u l=1u
M1271 n2480 net379 VSS VSS nmos w=1u l=1u
M1272 net379 n2414 net380 VSS nmos w=1u l=1u
M1273 net379 net377 net378 VSS nmos w=1u l=1u
M1274 net380 net378 VSS VSS nmos w=1u l=1u
M1275 net379 net377 net381 VDD pmos w=2u l=1u
M1276 net377 n2414 VDD VDD pmos w=2u l=1u
M1277 net378 n2414 net379 VDD pmos w=2u l=1u
M1278 net378 n2415 VDD VDD pmos w=2u l=1u
M1279 n2480 net379 VDD VDD pmos w=2u l=1u
M1280 net381 net378 VDD VDD pmos w=2u l=1u
M1281 n2415 n2486 VDD VDD pmos w=2u l=1u
M1282 n2415 n2486 VSS VSS nmos w=1u l=1u
M1283 n2479 n2488 net382 VSS nmos w=1u l=1u
M1284 net382 n2487 VSS VSS nmos w=1u l=1u
M1285 n2479 n2488 VDD VDD pmos w=2u l=1u
M1286 n2479 n2487 VDD VDD pmos w=2u l=1u
M1287 net383 n2486 VSS VSS nmos w=1u l=1u
M1288 net384 n2414 VSS VSS nmos w=1u l=1u
M1289 n2488 net385 VSS VSS nmos w=1u l=1u
M1290 net385 n2486 net386 VSS nmos w=1u l=1u
M1291 net385 net383 net384 VSS nmos w=1u l=1u
M1292 net386 net384 VSS VSS nmos w=1u l=1u
M1293 net385 net383 net387 VDD pmos w=2u l=1u
M1294 net383 n2486 VDD VDD pmos w=2u l=1u
M1295 net384 n2486 net385 VDD pmos w=2u l=1u
M1296 net384 n2414 VDD VDD pmos w=2u l=1u
M1297 n2488 net385 VDD VDD pmos w=2u l=1u
M1298 net387 net384 VDD VDD pmos w=2u l=1u
M1299 n2486 N494 net388 VSS nmos w=1u l=1u
M1300 net388 N188 VSS VSS nmos w=1u l=1u
M1301 n2486 N494 VDD VDD pmos w=2u l=1u
M1302 n2486 N188 VDD VDD pmos w=2u l=1u
M1303 n2414 n2413 net389 VSS nmos w=1u l=1u
M1304 net389 n2489 VSS VSS nmos w=1u l=1u
M1305 n2414 n2413 VDD VDD pmos w=2u l=1u
M1306 n2414 n2489 VDD VDD pmos w=2u l=1u
M1307 n2413 n2491 net390 VSS nmos w=1u l=1u
M1308 net390 n2490 VSS VSS nmos w=1u l=1u
M1309 n2413 n2491 VDD VDD pmos w=2u l=1u
M1310 n2413 n2490 VDD VDD pmos w=2u l=1u
M1311 n2491 n2493 net391 VSS nmos w=1u l=1u
M1312 net391 n2492 VSS VSS nmos w=1u l=1u
M1313 n2491 n2493 VDD VDD pmos w=2u l=1u
M1314 n2491 n2492 VDD VDD pmos w=2u l=1u
M1315 n2492 net392 VSS VSS nmos w=1u l=1u
M1316 net392 n2494 VSS VSS nmos w=1u l=1u
M1317 net392 n2495 VSS VSS nmos w=1u l=1u
M1318 net392 n2495 net393 VDD pmos w=2u l=1u
M1319 n2492 net392 VDD VDD pmos w=2u l=1u
M1320 net393 n2494 VDD VDD pmos w=2u l=1u
M1321 net394 n2424 VSS VSS nmos w=1u l=1u
M1322 net395 n2425 VSS VSS nmos w=1u l=1u
M1323 n2490 net396 VSS VSS nmos w=1u l=1u
M1324 net396 n2424 net397 VSS nmos w=1u l=1u
M1325 net396 net394 net395 VSS nmos w=1u l=1u
M1326 net397 net395 VSS VSS nmos w=1u l=1u
M1327 net396 net394 net398 VDD pmos w=2u l=1u
M1328 net394 n2424 VDD VDD pmos w=2u l=1u
M1329 net395 n2424 net396 VDD pmos w=2u l=1u
M1330 net395 n2425 VDD VDD pmos w=2u l=1u
M1331 n2490 net396 VDD VDD pmos w=2u l=1u
M1332 net398 net395 VDD VDD pmos w=2u l=1u
M1333 n2425 n2496 VDD VDD pmos w=2u l=1u
M1334 n2425 n2496 VSS VSS nmos w=1u l=1u
M1335 n2489 n2498 net399 VSS nmos w=1u l=1u
M1336 net399 n2497 VSS VSS nmos w=1u l=1u
M1337 n2489 n2498 VDD VDD pmos w=2u l=1u
M1338 n2489 n2497 VDD VDD pmos w=2u l=1u
M1339 net400 n2496 VSS VSS nmos w=1u l=1u
M1340 net401 n2424 VSS VSS nmos w=1u l=1u
M1341 n2498 net402 VSS VSS nmos w=1u l=1u
M1342 net402 n2496 net403 VSS nmos w=1u l=1u
M1343 net402 net400 net401 VSS nmos w=1u l=1u
M1344 net403 net401 VSS VSS nmos w=1u l=1u
M1345 net402 net400 net404 VDD pmos w=2u l=1u
M1346 net400 n2496 VDD VDD pmos w=2u l=1u
M1347 net401 n2496 net402 VDD pmos w=2u l=1u
M1348 net401 n2424 VDD VDD pmos w=2u l=1u
M1349 n2498 net402 VDD VDD pmos w=2u l=1u
M1350 net404 net401 VDD VDD pmos w=2u l=1u
M1351 n2496 N477 net405 VSS nmos w=1u l=1u
M1352 net405 N205 VSS VSS nmos w=1u l=1u
M1353 n2496 N477 VDD VDD pmos w=2u l=1u
M1354 n2496 N205 VDD VDD pmos w=2u l=1u
M1355 n2424 n2423 net406 VSS nmos w=1u l=1u
M1356 net406 n2499 VSS VSS nmos w=1u l=1u
M1357 n2424 n2423 VDD VDD pmos w=2u l=1u
M1358 n2424 n2499 VDD VDD pmos w=2u l=1u
M1359 n2423 n2501 net407 VSS nmos w=1u l=1u
M1360 net407 n2500 VSS VSS nmos w=1u l=1u
M1361 n2423 n2501 VDD VDD pmos w=2u l=1u
M1362 n2423 n2500 VDD VDD pmos w=2u l=1u
M1363 n2501 n2503 net408 VSS nmos w=1u l=1u
M1364 net408 n2502 VSS VSS nmos w=1u l=1u
M1365 n2501 n2503 VDD VDD pmos w=2u l=1u
M1366 n2501 n2502 VDD VDD pmos w=2u l=1u
M1367 n2502 n2505 net409 VSS nmos w=1u l=1u
M1368 net409 n2504 VSS VSS nmos w=1u l=1u
M1369 n2502 n2505 VDD VDD pmos w=2u l=1u
M1370 n2502 n2504 VDD VDD pmos w=2u l=1u
M1371 net410 n2435 VSS VSS nmos w=1u l=1u
M1372 net411 n2436 VSS VSS nmos w=1u l=1u
M1373 n2500 net412 VSS VSS nmos w=1u l=1u
M1374 net412 n2435 net413 VSS nmos w=1u l=1u
M1375 net412 net410 net411 VSS nmos w=1u l=1u
M1376 net413 net411 VSS VSS nmos w=1u l=1u
M1377 net412 net410 net414 VDD pmos w=2u l=1u
M1378 net410 n2435 VDD VDD pmos w=2u l=1u
M1379 net411 n2435 net412 VDD pmos w=2u l=1u
M1380 net411 n2436 VDD VDD pmos w=2u l=1u
M1381 n2500 net412 VDD VDD pmos w=2u l=1u
M1382 net414 net411 VDD VDD pmos w=2u l=1u
M1383 n2435 n2506 VDD VDD pmos w=2u l=1u
M1384 n2435 n2506 VSS VSS nmos w=1u l=1u
M1385 n2499 n2508 net415 VSS nmos w=1u l=1u
M1386 net415 n2507 VSS VSS nmos w=1u l=1u
M1387 n2499 n2508 VDD VDD pmos w=2u l=1u
M1388 n2499 n2507 VDD VDD pmos w=2u l=1u
M1389 net416 n2436 VSS VSS nmos w=1u l=1u
M1390 net417 n2506 VSS VSS nmos w=1u l=1u
M1391 n2508 net418 VSS VSS nmos w=1u l=1u
M1392 net418 n2436 net419 VSS nmos w=1u l=1u
M1393 net418 net416 net417 VSS nmos w=1u l=1u
M1394 net419 net417 VSS VSS nmos w=1u l=1u
M1395 net418 net416 net420 VDD pmos w=2u l=1u
M1396 net416 n2436 VDD VDD pmos w=2u l=1u
M1397 net417 n2436 net418 VDD pmos w=2u l=1u
M1398 net417 n2506 VDD VDD pmos w=2u l=1u
M1399 n2508 net418 VDD VDD pmos w=2u l=1u
M1400 net420 net417 VDD VDD pmos w=2u l=1u
M1401 n2436 N460 net421 VSS nmos w=1u l=1u
M1402 net421 N222 VSS VSS nmos w=1u l=1u
M1403 n2436 N460 VDD VDD pmos w=2u l=1u
M1404 n2436 N222 VDD VDD pmos w=2u l=1u
M1405 n2506 n2433 net422 VSS nmos w=1u l=1u
M1406 net422 n2509 VSS VSS nmos w=1u l=1u
M1407 n2506 n2433 VDD VDD pmos w=2u l=1u
M1408 n2506 n2509 VDD VDD pmos w=2u l=1u
M1409 n2433 n2511 net423 VSS nmos w=1u l=1u
M1410 net423 n2510 VSS VSS nmos w=1u l=1u
M1411 n2433 n2511 VDD VDD pmos w=2u l=1u
M1412 n2433 n2510 VDD VDD pmos w=2u l=1u
M1413 n2511 n2513 net424 VSS nmos w=1u l=1u
M1414 net424 n2512 VSS VSS nmos w=1u l=1u
M1415 n2511 n2513 VDD VDD pmos w=2u l=1u
M1416 n2511 n2512 VDD VDD pmos w=2u l=1u
M1417 n2509 n2512 net425 VSS nmos w=1u l=1u
M1418 net425 n2514 VSS VSS nmos w=1u l=1u
M1419 n2509 n2512 VDD VDD pmos w=2u l=1u
M1420 n2509 n2514 VDD VDD pmos w=2u l=1u
M1421 n2512 n2516 net426 VSS nmos w=1u l=1u
M1422 net426 n2515 VSS VSS nmos w=1u l=1u
M1423 n2512 n2516 VDD VDD pmos w=2u l=1u
M1424 n2512 n2515 VDD VDD pmos w=2u l=1u
M1425 n2514 n2510 VSS VSS nmos w=1u l=1u
M1426 n2514 n2517 VSS VSS nmos w=1u l=1u
M1427 n2514 n2510 net427 VDD pmos w=2u l=1u
M1428 net427 n2517 VDD VDD pmos w=2u l=1u
M1429 n2510 net428 VSS VSS nmos w=1u l=1u
M1430 net429 n2518 VSS VSS nmos w=1u l=1u
M1431 net428 n2448 net429 VSS nmos w=1u l=1u
M1432 net428 n2518 VDD VDD pmos w=2u l=1u
M1433 net428 n2448 VDD VDD pmos w=2u l=1u
M1434 n2510 net428 VDD VDD pmos w=2u l=1u
M1435 n2518 N443 net430 VSS nmos w=1u l=1u
M1436 net430 n2519 VSS VSS nmos w=1u l=1u
M1437 n2518 N443 VDD VDD pmos w=2u l=1u
M1438 n2518 n2519 VDD VDD pmos w=2u l=1u
M1439 n2519 n2521 VSS VSS nmos w=1u l=1u
M1440 n2519 n2520 VSS VSS nmos w=1u l=1u
M1441 n2519 n2521 net431 VDD pmos w=2u l=1u
M1442 net431 n2520 VDD VDD pmos w=2u l=1u
M1443 n2521 n2523 VSS VSS nmos w=1u l=1u
M1444 n2521 n2522 VSS VSS nmos w=1u l=1u
M1445 n2521 n2523 net432 VDD pmos w=2u l=1u
M1446 net432 n2522 VDD VDD pmos w=2u l=1u
M1447 n2523 n2270 net433 VSS nmos w=1u l=1u
M1448 net433 n2524 VSS VSS nmos w=1u l=1u
M1449 n2523 n2270 VDD VDD pmos w=2u l=1u
M1450 n2523 n2524 VDD VDD pmos w=2u l=1u
M1451 n2524 n2525 net434 VSS nmos w=1u l=1u
M1452 net434 N239 VSS VSS nmos w=1u l=1u
M1453 n2524 n2525 VDD VDD pmos w=2u l=1u
M1454 n2524 N239 VDD VDD pmos w=2u l=1u
M1455 n2522 n2451 VDD VDD pmos w=2u l=1u
M1456 n2522 n2451 VSS VSS nmos w=1u l=1u
M1457 n2520 n2451 VSS VSS nmos w=1u l=1u
M1458 n2520 N426 VSS VSS nmos w=1u l=1u
M1459 n2520 n2451 net435 VDD pmos w=2u l=1u
M1460 net435 N426 VDD VDD pmos w=2u l=1u
M1461 n2448 n2527 net436 VSS nmos w=1u l=1u
M1462 net436 n2526 VSS VSS nmos w=1u l=1u
M1463 n2448 n2527 VDD VDD pmos w=2u l=1u
M1464 n2448 n2526 VDD VDD pmos w=2u l=1u
M1465 n2527 N239 net437 VSS nmos w=1u l=1u
M1466 net437 N443 VSS VSS nmos w=1u l=1u
M1467 n2527 N239 VDD VDD pmos w=2u l=1u
M1468 n2527 N443 VDD VDD pmos w=2u l=1u
M1469 net438 n2450 VSS VSS nmos w=1u l=1u
M1470 net439 n2451 VSS VSS nmos w=1u l=1u
M1471 n2526 net440 VSS VSS nmos w=1u l=1u
M1472 net440 n2450 net441 VSS nmos w=1u l=1u
M1473 net440 net438 net439 VSS nmos w=1u l=1u
M1474 net441 net439 VSS VSS nmos w=1u l=1u
M1475 net440 net438 net442 VDD pmos w=2u l=1u
M1476 net438 n2450 VDD VDD pmos w=2u l=1u
M1477 net439 n2450 net440 VDD pmos w=2u l=1u
M1478 net439 n2451 VDD VDD pmos w=2u l=1u
M1479 n2526 net440 VDD VDD pmos w=2u l=1u
M1480 net442 net439 VDD VDD pmos w=2u l=1u
M1481 n2450 N256 net443 VSS nmos w=1u l=1u
M1482 net443 N426 VSS VSS nmos w=1u l=1u
M1483 n2450 N256 VDD VDD pmos w=2u l=1u
M1484 n2450 N426 VDD VDD pmos w=2u l=1u
M1485 n2451 n2529 net444 VSS nmos w=1u l=1u
M1486 net444 n2528 VSS VSS nmos w=1u l=1u
M1487 n2451 n2529 VDD VDD pmos w=2u l=1u
M1488 n2451 n2528 VDD VDD pmos w=2u l=1u
M1489 n2529 n2531 net445 VSS nmos w=1u l=1u
M1490 net445 n2530 VSS VSS nmos w=1u l=1u
M1491 n2529 n2531 VDD VDD pmos w=2u l=1u
M1492 n2529 n2530 VDD VDD pmos w=2u l=1u
M1493 n2517 n2513 VDD VDD pmos w=2u l=1u
M1494 n2517 n2513 VSS VSS nmos w=1u l=1u
M1495 n2507 n2533 VSS VSS nmos w=1u l=1u
M1496 n2507 n2532 VSS VSS nmos w=1u l=1u
M1497 n2507 n2533 net446 VDD pmos w=2u l=1u
M1498 net446 n2532 VDD VDD pmos w=2u l=1u
M1499 n2533 net447 VSS VSS nmos w=1u l=1u
M1500 net448 n2504 VSS VSS nmos w=1u l=1u
M1501 net447 n2505 net448 VSS nmos w=1u l=1u
M1502 net447 n2504 VDD VDD pmos w=2u l=1u
M1503 net447 n2505 VDD VDD pmos w=2u l=1u
M1504 n2533 net447 VDD VDD pmos w=2u l=1u
M1505 n2532 n2503 VDD VDD pmos w=2u l=1u
M1506 n2532 n2503 VSS VSS nmos w=1u l=1u
M1507 n2497 n2535 VSS VSS nmos w=1u l=1u
M1508 n2497 n2534 VSS VSS nmos w=1u l=1u
M1509 n2497 n2535 net449 VDD pmos w=2u l=1u
M1510 net449 n2534 VDD VDD pmos w=2u l=1u
M1511 n2535 n2494 VSS VSS nmos w=1u l=1u
M1512 n2535 n2495 VSS VSS nmos w=1u l=1u
M1513 n2535 n2494 net450 VDD pmos w=2u l=1u
M1514 net450 n2495 VDD VDD pmos w=2u l=1u
M1515 n2534 n2493 VDD VDD pmos w=2u l=1u
M1516 n2534 n2493 VSS VSS nmos w=1u l=1u
M1517 n2487 n2537 VSS VSS nmos w=1u l=1u
M1518 n2487 n2536 VSS VSS nmos w=1u l=1u
M1519 n2487 n2537 net451 VDD pmos w=2u l=1u
M1520 net451 n2536 VDD VDD pmos w=2u l=1u
M1521 n2537 n2484 VSS VSS nmos w=1u l=1u
M1522 n2537 n2485 VSS VSS nmos w=1u l=1u
M1523 n2537 n2484 net452 VDD pmos w=2u l=1u
M1524 net452 n2485 VDD VDD pmos w=2u l=1u
M1525 n2536 n2483 VDD VDD pmos w=2u l=1u
M1526 n2536 n2483 VSS VSS nmos w=1u l=1u
M1527 n2477 n2539 VSS VSS nmos w=1u l=1u
M1528 n2477 n2538 VSS VSS nmos w=1u l=1u
M1529 n2477 n2539 net453 VDD pmos w=2u l=1u
M1530 net453 n2538 VDD VDD pmos w=2u l=1u
M1531 n2539 n2474 VSS VSS nmos w=1u l=1u
M1532 n2539 n2475 VSS VSS nmos w=1u l=1u
M1533 n2539 n2474 net454 VDD pmos w=2u l=1u
M1534 net454 n2475 VDD VDD pmos w=2u l=1u
M1535 n2538 n2473 VDD VDD pmos w=2u l=1u
M1536 n2538 n2473 VSS VSS nmos w=1u l=1u
M1537 n2398 N528 net455 VSS nmos w=1u l=1u
M1538 net455 N154 VSS VSS nmos w=1u l=1u
M1539 n2398 N528 VDD VDD pmos w=2u l=1u
M1540 n2398 N154 VDD VDD pmos w=2u l=1u
M1541 N6220 n2540 net456 VSS nmos w=1u l=1u
M1542 net456 n2462 VSS VSS nmos w=1u l=1u
M1543 N6220 n2540 VDD VDD pmos w=2u l=1u
M1544 N6220 n2462 VDD VDD pmos w=2u l=1u
M1545 n2540 net457 VSS VSS nmos w=1u l=1u
M1546 net457 n2541 VSS VSS nmos w=1u l=1u
M1547 net457 n2542 VSS VSS nmos w=1u l=1u
M1548 net457 n2542 net458 VDD pmos w=2u l=1u
M1549 n2540 net457 VDD VDD pmos w=2u l=1u
M1550 net458 n2541 VDD VDD pmos w=2u l=1u
M1551 n2462 n2542 net459 VSS nmos w=1u l=1u
M1552 net459 n2541 VSS VSS nmos w=1u l=1u
M1553 n2462 n2542 VDD VDD pmos w=2u l=1u
M1554 n2462 n2541 VDD VDD pmos w=2u l=1u
M1555 n2542 n2544 net460 VSS nmos w=1u l=1u
M1556 net460 n2543 VSS VSS nmos w=1u l=1u
M1557 n2542 n2544 VDD VDD pmos w=2u l=1u
M1558 n2542 n2543 VDD VDD pmos w=2u l=1u
M1559 n2543 n2546 net461 VSS nmos w=1u l=1u
M1560 net461 n2545 VSS VSS nmos w=1u l=1u
M1561 n2543 n2546 VDD VDD pmos w=2u l=1u
M1562 n2543 n2545 VDD VDD pmos w=2u l=1u
M1563 net462 n2464 VSS VSS nmos w=1u l=1u
M1564 net463 n2463 VSS VSS nmos w=1u l=1u
M1565 n2541 net464 VSS VSS nmos w=1u l=1u
M1566 net464 n2464 net465 VSS nmos w=1u l=1u
M1567 net464 net462 net463 VSS nmos w=1u l=1u
M1568 net465 net463 VSS VSS nmos w=1u l=1u
M1569 net464 net462 net466 VDD pmos w=2u l=1u
M1570 net462 n2464 VDD VDD pmos w=2u l=1u
M1571 net463 n2464 net464 VDD pmos w=2u l=1u
M1572 net463 n2463 VDD VDD pmos w=2u l=1u
M1573 n2541 net464 VDD VDD pmos w=2u l=1u
M1574 net466 net463 VDD VDD pmos w=2u l=1u
M1575 n2464 n2548 net467 VSS nmos w=1u l=1u
M1576 net467 n2547 VSS VSS nmos w=1u l=1u
M1577 n2464 n2548 VDD VDD pmos w=2u l=1u
M1578 n2464 n2547 VDD VDD pmos w=2u l=1u
M1579 n2547 n2550 net468 VSS nmos w=1u l=1u
M1580 net468 n2549 VSS VSS nmos w=1u l=1u
M1581 n2547 n2550 VDD VDD pmos w=2u l=1u
M1582 n2547 n2549 VDD VDD pmos w=2u l=1u
M1583 net469 n2467 VSS VSS nmos w=1u l=1u
M1584 net470 n2468 VSS VSS nmos w=1u l=1u
M1585 n2463 net471 VSS VSS nmos w=1u l=1u
M1586 net471 n2467 net472 VSS nmos w=1u l=1u
M1587 net471 net469 net470 VSS nmos w=1u l=1u
M1588 net472 net470 VSS VSS nmos w=1u l=1u
M1589 net471 net469 net473 VDD pmos w=2u l=1u
M1590 net469 n2467 VDD VDD pmos w=2u l=1u
M1591 net470 n2467 net471 VDD pmos w=2u l=1u
M1592 net470 n2468 VDD VDD pmos w=2u l=1u
M1593 n2463 net471 VDD VDD pmos w=2u l=1u
M1594 net473 net470 VDD VDD pmos w=2u l=1u
M1595 n2467 net474 VSS VSS nmos w=1u l=1u
M1596 net475 n2466 VSS VSS nmos w=1u l=1u
M1597 net474 n2551 net475 VSS nmos w=1u l=1u
M1598 net474 n2466 VDD VDD pmos w=2u l=1u
M1599 net474 n2551 VDD VDD pmos w=2u l=1u
M1600 n2467 net474 VDD VDD pmos w=2u l=1u
M1601 n2466 n2553 net476 VSS nmos w=1u l=1u
M1602 net476 n2552 VSS VSS nmos w=1u l=1u
M1603 n2466 n2553 VDD VDD pmos w=2u l=1u
M1604 n2466 n2552 VDD VDD pmos w=2u l=1u
M1605 n2553 n2555 net477 VSS nmos w=1u l=1u
M1606 net477 n2554 VSS VSS nmos w=1u l=1u
M1607 n2553 n2555 VDD VDD pmos w=2u l=1u
M1608 n2553 n2554 VDD VDD pmos w=2u l=1u
M1609 n2554 net478 VSS VSS nmos w=1u l=1u
M1610 net478 n2556 VSS VSS nmos w=1u l=1u
M1611 net478 n2557 VSS VSS nmos w=1u l=1u
M1612 net478 n2557 net479 VDD pmos w=2u l=1u
M1613 n2554 net478 VDD VDD pmos w=2u l=1u
M1614 net479 n2556 VDD VDD pmos w=2u l=1u
M1615 net480 n2474 VSS VSS nmos w=1u l=1u
M1616 net481 n2475 VSS VSS nmos w=1u l=1u
M1617 n2552 net482 VSS VSS nmos w=1u l=1u
M1618 net482 n2474 net483 VSS nmos w=1u l=1u
M1619 net482 net480 net481 VSS nmos w=1u l=1u
M1620 net483 net481 VSS VSS nmos w=1u l=1u
M1621 net482 net480 net484 VDD pmos w=2u l=1u
M1622 net480 n2474 VDD VDD pmos w=2u l=1u
M1623 net481 n2474 net482 VDD pmos w=2u l=1u
M1624 net481 n2475 VDD VDD pmos w=2u l=1u
M1625 n2552 net482 VDD VDD pmos w=2u l=1u
M1626 net484 net481 VDD VDD pmos w=2u l=1u
M1627 n2475 n2558 VDD VDD pmos w=2u l=1u
M1628 n2475 n2558 VSS VSS nmos w=1u l=1u
M1629 n2551 n2560 net485 VSS nmos w=1u l=1u
M1630 net485 n2559 VSS VSS nmos w=1u l=1u
M1631 n2551 n2560 VDD VDD pmos w=2u l=1u
M1632 n2551 n2559 VDD VDD pmos w=2u l=1u
M1633 net486 n2558 VSS VSS nmos w=1u l=1u
M1634 net487 n2474 VSS VSS nmos w=1u l=1u
M1635 n2560 net488 VSS VSS nmos w=1u l=1u
M1636 net488 n2558 net489 VSS nmos w=1u l=1u
M1637 net488 net486 net487 VSS nmos w=1u l=1u
M1638 net489 net487 VSS VSS nmos w=1u l=1u
M1639 net488 net486 net490 VDD pmos w=2u l=1u
M1640 net486 n2558 VDD VDD pmos w=2u l=1u
M1641 net487 n2558 net488 VDD pmos w=2u l=1u
M1642 net487 n2474 VDD VDD pmos w=2u l=1u
M1643 n2560 net488 VDD VDD pmos w=2u l=1u
M1644 net490 net487 VDD VDD pmos w=2u l=1u
M1645 n2558 N511 net491 VSS nmos w=1u l=1u
M1646 net491 N154 VSS VSS nmos w=1u l=1u
M1647 n2558 N511 VDD VDD pmos w=2u l=1u
M1648 n2558 N154 VDD VDD pmos w=2u l=1u
M1649 n2474 n2473 net492 VSS nmos w=1u l=1u
M1650 net492 n2561 VSS VSS nmos w=1u l=1u
M1651 n2474 n2473 VDD VDD pmos w=2u l=1u
M1652 n2474 n2561 VDD VDD pmos w=2u l=1u
M1653 n2473 n2563 net493 VSS nmos w=1u l=1u
M1654 net493 n2562 VSS VSS nmos w=1u l=1u
M1655 n2473 n2563 VDD VDD pmos w=2u l=1u
M1656 n2473 n2562 VDD VDD pmos w=2u l=1u
M1657 n2563 n2565 net494 VSS nmos w=1u l=1u
M1658 net494 n2564 VSS VSS nmos w=1u l=1u
M1659 n2563 n2565 VDD VDD pmos w=2u l=1u
M1660 n2563 n2564 VDD VDD pmos w=2u l=1u
M1661 n2564 net495 VSS VSS nmos w=1u l=1u
M1662 net495 n2566 VSS VSS nmos w=1u l=1u
M1663 net495 n2567 VSS VSS nmos w=1u l=1u
M1664 net495 n2567 net496 VDD pmos w=2u l=1u
M1665 n2564 net495 VDD VDD pmos w=2u l=1u
M1666 net496 n2566 VDD VDD pmos w=2u l=1u
M1667 net497 n2484 VSS VSS nmos w=1u l=1u
M1668 net498 n2485 VSS VSS nmos w=1u l=1u
M1669 n2562 net499 VSS VSS nmos w=1u l=1u
M1670 net499 n2484 net500 VSS nmos w=1u l=1u
M1671 net499 net497 net498 VSS nmos w=1u l=1u
M1672 net500 net498 VSS VSS nmos w=1u l=1u
M1673 net499 net497 net501 VDD pmos w=2u l=1u
M1674 net497 n2484 VDD VDD pmos w=2u l=1u
M1675 net498 n2484 net499 VDD pmos w=2u l=1u
M1676 net498 n2485 VDD VDD pmos w=2u l=1u
M1677 n2562 net499 VDD VDD pmos w=2u l=1u
M1678 net501 net498 VDD VDD pmos w=2u l=1u
M1679 n2485 n2568 VDD VDD pmos w=2u l=1u
M1680 n2485 n2568 VSS VSS nmos w=1u l=1u
M1681 n2561 n2570 net502 VSS nmos w=1u l=1u
M1682 net502 n2569 VSS VSS nmos w=1u l=1u
M1683 n2561 n2570 VDD VDD pmos w=2u l=1u
M1684 n2561 n2569 VDD VDD pmos w=2u l=1u
M1685 net503 n2568 VSS VSS nmos w=1u l=1u
M1686 net504 n2484 VSS VSS nmos w=1u l=1u
M1687 n2570 net505 VSS VSS nmos w=1u l=1u
M1688 net505 n2568 net506 VSS nmos w=1u l=1u
M1689 net505 net503 net504 VSS nmos w=1u l=1u
M1690 net506 net504 VSS VSS nmos w=1u l=1u
M1691 net505 net503 net507 VDD pmos w=2u l=1u
M1692 net503 n2568 VDD VDD pmos w=2u l=1u
M1693 net504 n2568 net505 VDD pmos w=2u l=1u
M1694 net504 n2484 VDD VDD pmos w=2u l=1u
M1695 n2570 net505 VDD VDD pmos w=2u l=1u
M1696 net507 net504 VDD VDD pmos w=2u l=1u
M1697 n2568 N494 net508 VSS nmos w=1u l=1u
M1698 net508 N171 VSS VSS nmos w=1u l=1u
M1699 n2568 N494 VDD VDD pmos w=2u l=1u
M1700 n2568 N171 VDD VDD pmos w=2u l=1u
M1701 n2484 n2483 net509 VSS nmos w=1u l=1u
M1702 net509 n2571 VSS VSS nmos w=1u l=1u
M1703 n2484 n2483 VDD VDD pmos w=2u l=1u
M1704 n2484 n2571 VDD VDD pmos w=2u l=1u
M1705 n2483 n2573 net510 VSS nmos w=1u l=1u
M1706 net510 n2572 VSS VSS nmos w=1u l=1u
M1707 n2483 n2573 VDD VDD pmos w=2u l=1u
M1708 n2483 n2572 VDD VDD pmos w=2u l=1u
M1709 n2573 n2575 net511 VSS nmos w=1u l=1u
M1710 net511 n2574 VSS VSS nmos w=1u l=1u
M1711 n2573 n2575 VDD VDD pmos w=2u l=1u
M1712 n2573 n2574 VDD VDD pmos w=2u l=1u
M1713 n2574 net512 VSS VSS nmos w=1u l=1u
M1714 net512 n2576 VSS VSS nmos w=1u l=1u
M1715 net512 n2577 VSS VSS nmos w=1u l=1u
M1716 net512 n2577 net513 VDD pmos w=2u l=1u
M1717 n2574 net512 VDD VDD pmos w=2u l=1u
M1718 net513 n2576 VDD VDD pmos w=2u l=1u
M1719 net514 n2494 VSS VSS nmos w=1u l=1u
M1720 net515 n2495 VSS VSS nmos w=1u l=1u
M1721 n2572 net516 VSS VSS nmos w=1u l=1u
M1722 net516 n2494 net517 VSS nmos w=1u l=1u
M1723 net516 net514 net515 VSS nmos w=1u l=1u
M1724 net517 net515 VSS VSS nmos w=1u l=1u
M1725 net516 net514 net518 VDD pmos w=2u l=1u
M1726 net514 n2494 VDD VDD pmos w=2u l=1u
M1727 net515 n2494 net516 VDD pmos w=2u l=1u
M1728 net515 n2495 VDD VDD pmos w=2u l=1u
M1729 n2572 net516 VDD VDD pmos w=2u l=1u
M1730 net518 net515 VDD VDD pmos w=2u l=1u
M1731 n2495 n2578 VDD VDD pmos w=2u l=1u
M1732 n2495 n2578 VSS VSS nmos w=1u l=1u
M1733 n2571 n2580 net519 VSS nmos w=1u l=1u
M1734 net519 n2579 VSS VSS nmos w=1u l=1u
M1735 n2571 n2580 VDD VDD pmos w=2u l=1u
M1736 n2571 n2579 VDD VDD pmos w=2u l=1u
M1737 net520 n2578 VSS VSS nmos w=1u l=1u
M1738 net521 n2494 VSS VSS nmos w=1u l=1u
M1739 n2580 net522 VSS VSS nmos w=1u l=1u
M1740 net522 n2578 net523 VSS nmos w=1u l=1u
M1741 net522 net520 net521 VSS nmos w=1u l=1u
M1742 net523 net521 VSS VSS nmos w=1u l=1u
M1743 net522 net520 net524 VDD pmos w=2u l=1u
M1744 net520 n2578 VDD VDD pmos w=2u l=1u
M1745 net521 n2578 net522 VDD pmos w=2u l=1u
M1746 net521 n2494 VDD VDD pmos w=2u l=1u
M1747 n2580 net522 VDD VDD pmos w=2u l=1u
M1748 net524 net521 VDD VDD pmos w=2u l=1u
M1749 n2578 N477 net525 VSS nmos w=1u l=1u
M1750 net525 N188 VSS VSS nmos w=1u l=1u
M1751 n2578 N477 VDD VDD pmos w=2u l=1u
M1752 n2578 N188 VDD VDD pmos w=2u l=1u
M1753 n2494 n2493 net526 VSS nmos w=1u l=1u
M1754 net526 n2581 VSS VSS nmos w=1u l=1u
M1755 n2494 n2493 VDD VDD pmos w=2u l=1u
M1756 n2494 n2581 VDD VDD pmos w=2u l=1u
M1757 n2493 n2583 net527 VSS nmos w=1u l=1u
M1758 net527 n2582 VSS VSS nmos w=1u l=1u
M1759 n2493 n2583 VDD VDD pmos w=2u l=1u
M1760 n2493 n2582 VDD VDD pmos w=2u l=1u
M1761 n2583 n2585 net528 VSS nmos w=1u l=1u
M1762 net528 n2584 VSS VSS nmos w=1u l=1u
M1763 n2583 n2585 VDD VDD pmos w=2u l=1u
M1764 n2583 n2584 VDD VDD pmos w=2u l=1u
M1765 n2584 net529 VSS VSS nmos w=1u l=1u
M1766 net529 n2586 VSS VSS nmos w=1u l=1u
M1767 net529 n2587 VSS VSS nmos w=1u l=1u
M1768 net529 n2587 net530 VDD pmos w=2u l=1u
M1769 n2584 net529 VDD VDD pmos w=2u l=1u
M1770 net530 n2586 VDD VDD pmos w=2u l=1u
M1771 net531 n2504 VSS VSS nmos w=1u l=1u
M1772 net532 n2505 VSS VSS nmos w=1u l=1u
M1773 n2582 net533 VSS VSS nmos w=1u l=1u
M1774 net533 n2504 net534 VSS nmos w=1u l=1u
M1775 net533 net531 net532 VSS nmos w=1u l=1u
M1776 net534 net532 VSS VSS nmos w=1u l=1u
M1777 net533 net531 net535 VDD pmos w=2u l=1u
M1778 net531 n2504 VDD VDD pmos w=2u l=1u
M1779 net532 n2504 net533 VDD pmos w=2u l=1u
M1780 net532 n2505 VDD VDD pmos w=2u l=1u
M1781 n2582 net533 VDD VDD pmos w=2u l=1u
M1782 net535 net532 VDD VDD pmos w=2u l=1u
M1783 n2504 n2588 VDD VDD pmos w=2u l=1u
M1784 n2504 n2588 VSS VSS nmos w=1u l=1u
M1785 n2581 n2590 net536 VSS nmos w=1u l=1u
M1786 net536 n2589 VSS VSS nmos w=1u l=1u
M1787 n2581 n2590 VDD VDD pmos w=2u l=1u
M1788 n2581 n2589 VDD VDD pmos w=2u l=1u
M1789 net537 n2505 VSS VSS nmos w=1u l=1u
M1790 net538 n2588 VSS VSS nmos w=1u l=1u
M1791 n2590 net539 VSS VSS nmos w=1u l=1u
M1792 net539 n2505 net540 VSS nmos w=1u l=1u
M1793 net539 net537 net538 VSS nmos w=1u l=1u
M1794 net540 net538 VSS VSS nmos w=1u l=1u
M1795 net539 net537 net541 VDD pmos w=2u l=1u
M1796 net537 n2505 VDD VDD pmos w=2u l=1u
M1797 net538 n2505 net539 VDD pmos w=2u l=1u
M1798 net538 n2588 VDD VDD pmos w=2u l=1u
M1799 n2590 net539 VDD VDD pmos w=2u l=1u
M1800 net541 net538 VDD VDD pmos w=2u l=1u
M1801 n2505 N460 net542 VSS nmos w=1u l=1u
M1802 net542 N205 VSS VSS nmos w=1u l=1u
M1803 n2505 N460 VDD VDD pmos w=2u l=1u
M1804 n2505 N205 VDD VDD pmos w=2u l=1u
M1805 n2588 n2503 net543 VSS nmos w=1u l=1u
M1806 net543 n2591 VSS VSS nmos w=1u l=1u
M1807 n2588 n2503 VDD VDD pmos w=2u l=1u
M1808 n2588 n2591 VDD VDD pmos w=2u l=1u
M1809 n2503 n2593 net544 VSS nmos w=1u l=1u
M1810 net544 n2592 VSS VSS nmos w=1u l=1u
M1811 n2503 n2593 VDD VDD pmos w=2u l=1u
M1812 n2503 n2592 VDD VDD pmos w=2u l=1u
M1813 n2593 n2595 net545 VSS nmos w=1u l=1u
M1814 net545 n2594 VSS VSS nmos w=1u l=1u
M1815 n2593 n2595 VDD VDD pmos w=2u l=1u
M1816 n2593 n2594 VDD VDD pmos w=2u l=1u
M1817 n2594 net546 VSS VSS nmos w=1u l=1u
M1818 net546 n2596 VSS VSS nmos w=1u l=1u
M1819 net546 n2597 VSS VSS nmos w=1u l=1u
M1820 net546 n2597 net547 VDD pmos w=2u l=1u
M1821 n2594 net546 VDD VDD pmos w=2u l=1u
M1822 net547 n2596 VDD VDD pmos w=2u l=1u
M1823 net548 n2515 VSS VSS nmos w=1u l=1u
M1824 net549 n2516 VSS VSS nmos w=1u l=1u
M1825 n2592 net550 VSS VSS nmos w=1u l=1u
M1826 net550 n2515 net551 VSS nmos w=1u l=1u
M1827 net550 net548 net549 VSS nmos w=1u l=1u
M1828 net551 net549 VSS VSS nmos w=1u l=1u
M1829 net550 net548 net552 VDD pmos w=2u l=1u
M1830 net548 n2515 VDD VDD pmos w=2u l=1u
M1831 net549 n2515 net550 VDD pmos w=2u l=1u
M1832 net549 n2516 VDD VDD pmos w=2u l=1u
M1833 n2592 net550 VDD VDD pmos w=2u l=1u
M1834 net552 net549 VDD VDD pmos w=2u l=1u
M1835 n2515 n2598 VDD VDD pmos w=2u l=1u
M1836 n2515 n2598 VSS VSS nmos w=1u l=1u
M1837 n2591 n2600 net553 VSS nmos w=1u l=1u
M1838 net553 n2599 VSS VSS nmos w=1u l=1u
M1839 n2591 n2600 VDD VDD pmos w=2u l=1u
M1840 n2591 n2599 VDD VDD pmos w=2u l=1u
M1841 net554 n2516 VSS VSS nmos w=1u l=1u
M1842 net555 n2598 VSS VSS nmos w=1u l=1u
M1843 n2600 net556 VSS VSS nmos w=1u l=1u
M1844 net556 n2516 net557 VSS nmos w=1u l=1u
M1845 net556 net554 net555 VSS nmos w=1u l=1u
M1846 net557 net555 VSS VSS nmos w=1u l=1u
M1847 net556 net554 net558 VDD pmos w=2u l=1u
M1848 net554 n2516 VDD VDD pmos w=2u l=1u
M1849 net555 n2516 net556 VDD pmos w=2u l=1u
M1850 net555 n2598 VDD VDD pmos w=2u l=1u
M1851 n2600 net556 VDD VDD pmos w=2u l=1u
M1852 net558 net555 VDD VDD pmos w=2u l=1u
M1853 n2516 N443 net559 VSS nmos w=1u l=1u
M1854 net559 N222 VSS VSS nmos w=1u l=1u
M1855 n2516 N443 VDD VDD pmos w=2u l=1u
M1856 n2516 N222 VDD VDD pmos w=2u l=1u
M1857 n2598 n2513 net560 VSS nmos w=1u l=1u
M1858 net560 n2601 VSS VSS nmos w=1u l=1u
M1859 n2598 n2513 VDD VDD pmos w=2u l=1u
M1860 n2598 n2601 VDD VDD pmos w=2u l=1u
M1861 n2513 n2603 net561 VSS nmos w=1u l=1u
M1862 net561 n2602 VSS VSS nmos w=1u l=1u
M1863 n2513 n2603 VDD VDD pmos w=2u l=1u
M1864 n2513 n2602 VDD VDD pmos w=2u l=1u
M1865 n2603 n2605 net562 VSS nmos w=1u l=1u
M1866 net562 n2604 VSS VSS nmos w=1u l=1u
M1867 n2603 n2605 VDD VDD pmos w=2u l=1u
M1868 n2603 n2604 VDD VDD pmos w=2u l=1u
M1869 n2601 n2604 net563 VSS nmos w=1u l=1u
M1870 net563 n2606 VSS VSS nmos w=1u l=1u
M1871 n2601 n2604 VDD VDD pmos w=2u l=1u
M1872 n2601 n2606 VDD VDD pmos w=2u l=1u
M1873 n2604 n2608 net564 VSS nmos w=1u l=1u
M1874 net564 n2607 VSS VSS nmos w=1u l=1u
M1875 n2604 n2608 VDD VDD pmos w=2u l=1u
M1876 n2604 n2607 VDD VDD pmos w=2u l=1u
M1877 n2606 n2602 VSS VSS nmos w=1u l=1u
M1878 n2606 n2609 VSS VSS nmos w=1u l=1u
M1879 n2606 n2602 net565 VDD pmos w=2u l=1u
M1880 net565 n2609 VDD VDD pmos w=2u l=1u
M1881 n2602 net566 VSS VSS nmos w=1u l=1u
M1882 net567 n2610 VSS VSS nmos w=1u l=1u
M1883 net566 n2528 net567 VSS nmos w=1u l=1u
M1884 net566 n2610 VDD VDD pmos w=2u l=1u
M1885 net566 n2528 VDD VDD pmos w=2u l=1u
M1886 n2602 net566 VDD VDD pmos w=2u l=1u
M1887 n2610 N426 net568 VSS nmos w=1u l=1u
M1888 net568 n2611 VSS VSS nmos w=1u l=1u
M1889 n2610 N426 VDD VDD pmos w=2u l=1u
M1890 n2610 n2611 VDD VDD pmos w=2u l=1u
M1891 n2611 n2613 VSS VSS nmos w=1u l=1u
M1892 n2611 n2612 VSS VSS nmos w=1u l=1u
M1893 n2611 n2613 net569 VDD pmos w=2u l=1u
M1894 net569 n2612 VDD VDD pmos w=2u l=1u
M1895 n2613 n2615 VSS VSS nmos w=1u l=1u
M1896 n2613 n2614 VSS VSS nmos w=1u l=1u
M1897 n2613 n2615 net570 VDD pmos w=2u l=1u
M1898 net570 n2614 VDD VDD pmos w=2u l=1u
M1899 n2615 n2270 net571 VSS nmos w=1u l=1u
M1900 net571 n2616 VSS VSS nmos w=1u l=1u
M1901 n2615 n2270 VDD VDD pmos w=2u l=1u
M1902 n2615 n2616 VDD VDD pmos w=2u l=1u
M1903 n2616 n2617 net572 VSS nmos w=1u l=1u
M1904 net572 N239 VSS VSS nmos w=1u l=1u
M1905 n2616 n2617 VDD VDD pmos w=2u l=1u
M1906 n2616 N239 VDD VDD pmos w=2u l=1u
M1907 n2614 n2531 VDD VDD pmos w=2u l=1u
M1908 n2614 n2531 VSS VSS nmos w=1u l=1u
M1909 n2612 n2531 VSS VSS nmos w=1u l=1u
M1910 n2612 N409 VSS VSS nmos w=1u l=1u
M1911 n2612 n2531 net573 VDD pmos w=2u l=1u
M1912 net573 N409 VDD VDD pmos w=2u l=1u
M1913 n2528 n2619 net574 VSS nmos w=1u l=1u
M1914 net574 n2618 VSS VSS nmos w=1u l=1u
M1915 n2528 n2619 VDD VDD pmos w=2u l=1u
M1916 n2528 n2618 VDD VDD pmos w=2u l=1u
M1917 n2619 N239 net575 VSS nmos w=1u l=1u
M1918 net575 N426 VSS VSS nmos w=1u l=1u
M1919 n2619 N239 VDD VDD pmos w=2u l=1u
M1920 n2619 N426 VDD VDD pmos w=2u l=1u
M1921 net576 n2530 VSS VSS nmos w=1u l=1u
M1922 net577 n2531 VSS VSS nmos w=1u l=1u
M1923 n2618 net578 VSS VSS nmos w=1u l=1u
M1924 net578 n2530 net579 VSS nmos w=1u l=1u
M1925 net578 net576 net577 VSS nmos w=1u l=1u
M1926 net579 net577 VSS VSS nmos w=1u l=1u
M1927 net578 net576 net580 VDD pmos w=2u l=1u
M1928 net576 n2530 VDD VDD pmos w=2u l=1u
M1929 net577 n2530 net578 VDD pmos w=2u l=1u
M1930 net577 n2531 VDD VDD pmos w=2u l=1u
M1931 n2618 net578 VDD VDD pmos w=2u l=1u
M1932 net580 net577 VDD VDD pmos w=2u l=1u
M1933 n2530 N256 net581 VSS nmos w=1u l=1u
M1934 net581 N409 VSS VSS nmos w=1u l=1u
M1935 n2530 N256 VDD VDD pmos w=2u l=1u
M1936 n2530 N409 VDD VDD pmos w=2u l=1u
M1937 n2531 n2621 net582 VSS nmos w=1u l=1u
M1938 net582 n2620 VSS VSS nmos w=1u l=1u
M1939 n2531 n2621 VDD VDD pmos w=2u l=1u
M1940 n2531 n2620 VDD VDD pmos w=2u l=1u
M1941 n2621 n2623 net583 VSS nmos w=1u l=1u
M1942 net583 n2622 VSS VSS nmos w=1u l=1u
M1943 n2621 n2623 VDD VDD pmos w=2u l=1u
M1944 n2621 n2622 VDD VDD pmos w=2u l=1u
M1945 n2609 n2605 VDD VDD pmos w=2u l=1u
M1946 n2609 n2605 VSS VSS nmos w=1u l=1u
M1947 n2599 n2625 VSS VSS nmos w=1u l=1u
M1948 n2599 n2624 VSS VSS nmos w=1u l=1u
M1949 n2599 n2625 net584 VDD pmos w=2u l=1u
M1950 net584 n2624 VDD VDD pmos w=2u l=1u
M1951 n2625 n2596 VSS VSS nmos w=1u l=1u
M1952 n2625 n2597 VSS VSS nmos w=1u l=1u
M1953 n2625 n2596 net585 VDD pmos w=2u l=1u
M1954 net585 n2597 VDD VDD pmos w=2u l=1u
M1955 n2624 n2595 VDD VDD pmos w=2u l=1u
M1956 n2624 n2595 VSS VSS nmos w=1u l=1u
M1957 n2589 n2627 VSS VSS nmos w=1u l=1u
M1958 n2589 n2626 VSS VSS nmos w=1u l=1u
M1959 n2589 n2627 net586 VDD pmos w=2u l=1u
M1960 net586 n2626 VDD VDD pmos w=2u l=1u
M1961 n2627 n2586 VSS VSS nmos w=1u l=1u
M1962 n2627 n2587 VSS VSS nmos w=1u l=1u
M1963 n2627 n2586 net587 VDD pmos w=2u l=1u
M1964 net587 n2587 VDD VDD pmos w=2u l=1u
M1965 n2626 n2585 VDD VDD pmos w=2u l=1u
M1966 n2626 n2585 VSS VSS nmos w=1u l=1u
M1967 n2579 n2629 VSS VSS nmos w=1u l=1u
M1968 n2579 n2628 VSS VSS nmos w=1u l=1u
M1969 n2579 n2629 net588 VDD pmos w=2u l=1u
M1970 net588 n2628 VDD VDD pmos w=2u l=1u
M1971 n2629 n2576 VSS VSS nmos w=1u l=1u
M1972 n2629 n2577 VSS VSS nmos w=1u l=1u
M1973 n2629 n2576 net589 VDD pmos w=2u l=1u
M1974 net589 n2577 VDD VDD pmos w=2u l=1u
M1975 n2628 n2575 VDD VDD pmos w=2u l=1u
M1976 n2628 n2575 VSS VSS nmos w=1u l=1u
M1977 n2569 n2631 VSS VSS nmos w=1u l=1u
M1978 n2569 n2630 VSS VSS nmos w=1u l=1u
M1979 n2569 n2631 net590 VDD pmos w=2u l=1u
M1980 net590 n2630 VDD VDD pmos w=2u l=1u
M1981 n2631 n2566 VSS VSS nmos w=1u l=1u
M1982 n2631 n2567 VSS VSS nmos w=1u l=1u
M1983 n2631 n2566 net591 VDD pmos w=2u l=1u
M1984 net591 n2567 VDD VDD pmos w=2u l=1u
M1985 n2630 n2565 VDD VDD pmos w=2u l=1u
M1986 n2630 n2565 VSS VSS nmos w=1u l=1u
M1987 n2559 n2633 VSS VSS nmos w=1u l=1u
M1988 n2559 n2632 VSS VSS nmos w=1u l=1u
M1989 n2559 n2633 net592 VDD pmos w=2u l=1u
M1990 net592 n2632 VDD VDD pmos w=2u l=1u
M1991 n2633 n2556 VSS VSS nmos w=1u l=1u
M1992 n2633 n2557 VSS VSS nmos w=1u l=1u
M1993 n2633 n2556 net593 VDD pmos w=2u l=1u
M1994 net593 n2557 VDD VDD pmos w=2u l=1u
M1995 n2632 n2555 VDD VDD pmos w=2u l=1u
M1996 n2632 n2555 VSS VSS nmos w=1u l=1u
M1997 n2468 N528 net594 VSS nmos w=1u l=1u
M1998 net594 N137 VSS VSS nmos w=1u l=1u
M1999 n2468 N528 VDD VDD pmos w=2u l=1u
M2000 n2468 N137 VDD VDD pmos w=2u l=1u
M2001 N6210 n2634 net595 VSS nmos w=1u l=1u
M2002 net595 n2544 VSS VSS nmos w=1u l=1u
M2003 N6210 n2634 VDD VDD pmos w=2u l=1u
M2004 N6210 n2544 VDD VDD pmos w=2u l=1u
M2005 n2634 net596 VSS VSS nmos w=1u l=1u
M2006 net596 n2635 VSS VSS nmos w=1u l=1u
M2007 net596 n2636 VSS VSS nmos w=1u l=1u
M2008 net596 n2636 net597 VDD pmos w=2u l=1u
M2009 n2634 net596 VDD VDD pmos w=2u l=1u
M2010 net597 n2635 VDD VDD pmos w=2u l=1u
M2011 n2544 n2636 net598 VSS nmos w=1u l=1u
M2012 net598 n2635 VSS VSS nmos w=1u l=1u
M2013 n2544 n2636 VDD VDD pmos w=2u l=1u
M2014 n2544 n2635 VDD VDD pmos w=2u l=1u
M2015 n2636 n2638 net599 VSS nmos w=1u l=1u
M2016 net599 n2637 VSS VSS nmos w=1u l=1u
M2017 n2636 n2638 VDD VDD pmos w=2u l=1u
M2018 n2636 n2637 VDD VDD pmos w=2u l=1u
M2019 n2637 n2640 net600 VSS nmos w=1u l=1u
M2020 net600 n2639 VSS VSS nmos w=1u l=1u
M2021 n2637 n2640 VDD VDD pmos w=2u l=1u
M2022 n2637 n2639 VDD VDD pmos w=2u l=1u
M2023 net601 n2546 VSS VSS nmos w=1u l=1u
M2024 net602 n2545 VSS VSS nmos w=1u l=1u
M2025 n2635 net603 VSS VSS nmos w=1u l=1u
M2026 net603 n2546 net604 VSS nmos w=1u l=1u
M2027 net603 net601 net602 VSS nmos w=1u l=1u
M2028 net604 net602 VSS VSS nmos w=1u l=1u
M2029 net603 net601 net605 VDD pmos w=2u l=1u
M2030 net601 n2546 VDD VDD pmos w=2u l=1u
M2031 net602 n2546 net603 VDD pmos w=2u l=1u
M2032 net602 n2545 VDD VDD pmos w=2u l=1u
M2033 n2635 net603 VDD VDD pmos w=2u l=1u
M2034 net605 net602 VDD VDD pmos w=2u l=1u
M2035 n2546 n2642 net606 VSS nmos w=1u l=1u
M2036 net606 n2641 VSS VSS nmos w=1u l=1u
M2037 n2546 n2642 VDD VDD pmos w=2u l=1u
M2038 n2546 n2641 VDD VDD pmos w=2u l=1u
M2039 n2641 n2644 net607 VSS nmos w=1u l=1u
M2040 net607 n2643 VSS VSS nmos w=1u l=1u
M2041 n2641 n2644 VDD VDD pmos w=2u l=1u
M2042 n2641 n2643 VDD VDD pmos w=2u l=1u
M2043 net608 n2549 VSS VSS nmos w=1u l=1u
M2044 net609 n2550 VSS VSS nmos w=1u l=1u
M2045 n2545 net610 VSS VSS nmos w=1u l=1u
M2046 net610 n2549 net611 VSS nmos w=1u l=1u
M2047 net610 net608 net609 VSS nmos w=1u l=1u
M2048 net611 net609 VSS VSS nmos w=1u l=1u
M2049 net610 net608 net612 VDD pmos w=2u l=1u
M2050 net608 n2549 VDD VDD pmos w=2u l=1u
M2051 net609 n2549 net610 VDD pmos w=2u l=1u
M2052 net609 n2550 VDD VDD pmos w=2u l=1u
M2053 n2545 net610 VDD VDD pmos w=2u l=1u
M2054 net612 net609 VDD VDD pmos w=2u l=1u
M2055 n2549 net613 VSS VSS nmos w=1u l=1u
M2056 net614 n2548 VSS VSS nmos w=1u l=1u
M2057 net613 n2645 net614 VSS nmos w=1u l=1u
M2058 net613 n2548 VDD VDD pmos w=2u l=1u
M2059 net613 n2645 VDD VDD pmos w=2u l=1u
M2060 n2549 net613 VDD VDD pmos w=2u l=1u
M2061 n2548 n2647 net615 VSS nmos w=1u l=1u
M2062 net615 n2646 VSS VSS nmos w=1u l=1u
M2063 n2548 n2647 VDD VDD pmos w=2u l=1u
M2064 n2548 n2646 VDD VDD pmos w=2u l=1u
M2065 n2647 n2649 net616 VSS nmos w=1u l=1u
M2066 net616 n2648 VSS VSS nmos w=1u l=1u
M2067 n2647 n2649 VDD VDD pmos w=2u l=1u
M2068 n2647 n2648 VDD VDD pmos w=2u l=1u
M2069 n2648 net617 VSS VSS nmos w=1u l=1u
M2070 net617 n2650 VSS VSS nmos w=1u l=1u
M2071 net617 n2651 VSS VSS nmos w=1u l=1u
M2072 net617 n2651 net618 VDD pmos w=2u l=1u
M2073 n2648 net617 VDD VDD pmos w=2u l=1u
M2074 net618 n2650 VDD VDD pmos w=2u l=1u
M2075 net619 n2556 VSS VSS nmos w=1u l=1u
M2076 net620 n2557 VSS VSS nmos w=1u l=1u
M2077 n2646 net621 VSS VSS nmos w=1u l=1u
M2078 net621 n2556 net622 VSS nmos w=1u l=1u
M2079 net621 net619 net620 VSS nmos w=1u l=1u
M2080 net622 net620 VSS VSS nmos w=1u l=1u
M2081 net621 net619 net623 VDD pmos w=2u l=1u
M2082 net619 n2556 VDD VDD pmos w=2u l=1u
M2083 net620 n2556 net621 VDD pmos w=2u l=1u
M2084 net620 n2557 VDD VDD pmos w=2u l=1u
M2085 n2646 net621 VDD VDD pmos w=2u l=1u
M2086 net623 net620 VDD VDD pmos w=2u l=1u
M2087 n2557 n2652 VDD VDD pmos w=2u l=1u
M2088 n2557 n2652 VSS VSS nmos w=1u l=1u
M2089 n2645 n2654 net624 VSS nmos w=1u l=1u
M2090 net624 n2653 VSS VSS nmos w=1u l=1u
M2091 n2645 n2654 VDD VDD pmos w=2u l=1u
M2092 n2645 n2653 VDD VDD pmos w=2u l=1u
M2093 net625 n2652 VSS VSS nmos w=1u l=1u
M2094 net626 n2556 VSS VSS nmos w=1u l=1u
M2095 n2654 net627 VSS VSS nmos w=1u l=1u
M2096 net627 n2652 net628 VSS nmos w=1u l=1u
M2097 net627 net625 net626 VSS nmos w=1u l=1u
M2098 net628 net626 VSS VSS nmos w=1u l=1u
M2099 net627 net625 net629 VDD pmos w=2u l=1u
M2100 net625 n2652 VDD VDD pmos w=2u l=1u
M2101 net626 n2652 net627 VDD pmos w=2u l=1u
M2102 net626 n2556 VDD VDD pmos w=2u l=1u
M2103 n2654 net627 VDD VDD pmos w=2u l=1u
M2104 net629 net626 VDD VDD pmos w=2u l=1u
M2105 n2652 N511 net630 VSS nmos w=1u l=1u
M2106 net630 N137 VSS VSS nmos w=1u l=1u
M2107 n2652 N511 VDD VDD pmos w=2u l=1u
M2108 n2652 N137 VDD VDD pmos w=2u l=1u
M2109 n2556 n2555 net631 VSS nmos w=1u l=1u
M2110 net631 n2655 VSS VSS nmos w=1u l=1u
M2111 n2556 n2555 VDD VDD pmos w=2u l=1u
M2112 n2556 n2655 VDD VDD pmos w=2u l=1u
M2113 n2555 n2657 net632 VSS nmos w=1u l=1u
M2114 net632 n2656 VSS VSS nmos w=1u l=1u
M2115 n2555 n2657 VDD VDD pmos w=2u l=1u
M2116 n2555 n2656 VDD VDD pmos w=2u l=1u
M2117 n2657 n2659 net633 VSS nmos w=1u l=1u
M2118 net633 n2658 VSS VSS nmos w=1u l=1u
M2119 n2657 n2659 VDD VDD pmos w=2u l=1u
M2120 n2657 n2658 VDD VDD pmos w=2u l=1u
M2121 n2658 net634 VSS VSS nmos w=1u l=1u
M2122 net634 n2660 VSS VSS nmos w=1u l=1u
M2123 net634 n2661 VSS VSS nmos w=1u l=1u
M2124 net634 n2661 net635 VDD pmos w=2u l=1u
M2125 n2658 net634 VDD VDD pmos w=2u l=1u
M2126 net635 n2660 VDD VDD pmos w=2u l=1u
M2127 net636 n2566 VSS VSS nmos w=1u l=1u
M2128 net637 n2567 VSS VSS nmos w=1u l=1u
M2129 n2656 net638 VSS VSS nmos w=1u l=1u
M2130 net638 n2566 net639 VSS nmos w=1u l=1u
M2131 net638 net636 net637 VSS nmos w=1u l=1u
M2132 net639 net637 VSS VSS nmos w=1u l=1u
M2133 net638 net636 net640 VDD pmos w=2u l=1u
M2134 net636 n2566 VDD VDD pmos w=2u l=1u
M2135 net637 n2566 net638 VDD pmos w=2u l=1u
M2136 net637 n2567 VDD VDD pmos w=2u l=1u
M2137 n2656 net638 VDD VDD pmos w=2u l=1u
M2138 net640 net637 VDD VDD pmos w=2u l=1u
M2139 n2567 n2662 VDD VDD pmos w=2u l=1u
M2140 n2567 n2662 VSS VSS nmos w=1u l=1u
M2141 n2655 n2664 net641 VSS nmos w=1u l=1u
M2142 net641 n2663 VSS VSS nmos w=1u l=1u
M2143 n2655 n2664 VDD VDD pmos w=2u l=1u
M2144 n2655 n2663 VDD VDD pmos w=2u l=1u
M2145 net642 n2662 VSS VSS nmos w=1u l=1u
M2146 net643 n2566 VSS VSS nmos w=1u l=1u
M2147 n2664 net644 VSS VSS nmos w=1u l=1u
M2148 net644 n2662 net645 VSS nmos w=1u l=1u
M2149 net644 net642 net643 VSS nmos w=1u l=1u
M2150 net645 net643 VSS VSS nmos w=1u l=1u
M2151 net644 net642 net646 VDD pmos w=2u l=1u
M2152 net642 n2662 VDD VDD pmos w=2u l=1u
M2153 net643 n2662 net644 VDD pmos w=2u l=1u
M2154 net643 n2566 VDD VDD pmos w=2u l=1u
M2155 n2664 net644 VDD VDD pmos w=2u l=1u
M2156 net646 net643 VDD VDD pmos w=2u l=1u
M2157 n2662 N494 net647 VSS nmos w=1u l=1u
M2158 net647 N154 VSS VSS nmos w=1u l=1u
M2159 n2662 N494 VDD VDD pmos w=2u l=1u
M2160 n2662 N154 VDD VDD pmos w=2u l=1u
M2161 n2566 n2565 net648 VSS nmos w=1u l=1u
M2162 net648 n2665 VSS VSS nmos w=1u l=1u
M2163 n2566 n2565 VDD VDD pmos w=2u l=1u
M2164 n2566 n2665 VDD VDD pmos w=2u l=1u
M2165 n2565 n2667 net649 VSS nmos w=1u l=1u
M2166 net649 n2666 VSS VSS nmos w=1u l=1u
M2167 n2565 n2667 VDD VDD pmos w=2u l=1u
M2168 n2565 n2666 VDD VDD pmos w=2u l=1u
M2169 n2667 n2669 net650 VSS nmos w=1u l=1u
M2170 net650 n2668 VSS VSS nmos w=1u l=1u
M2171 n2667 n2669 VDD VDD pmos w=2u l=1u
M2172 n2667 n2668 VDD VDD pmos w=2u l=1u
M2173 n2668 net651 VSS VSS nmos w=1u l=1u
M2174 net651 n2670 VSS VSS nmos w=1u l=1u
M2175 net651 n2671 VSS VSS nmos w=1u l=1u
M2176 net651 n2671 net652 VDD pmos w=2u l=1u
M2177 n2668 net651 VDD VDD pmos w=2u l=1u
M2178 net652 n2670 VDD VDD pmos w=2u l=1u
M2179 net653 n2576 VSS VSS nmos w=1u l=1u
M2180 net654 n2577 VSS VSS nmos w=1u l=1u
M2181 n2666 net655 VSS VSS nmos w=1u l=1u
M2182 net655 n2576 net656 VSS nmos w=1u l=1u
M2183 net655 net653 net654 VSS nmos w=1u l=1u
M2184 net656 net654 VSS VSS nmos w=1u l=1u
M2185 net655 net653 net657 VDD pmos w=2u l=1u
M2186 net653 n2576 VDD VDD pmos w=2u l=1u
M2187 net654 n2576 net655 VDD pmos w=2u l=1u
M2188 net654 n2577 VDD VDD pmos w=2u l=1u
M2189 n2666 net655 VDD VDD pmos w=2u l=1u
M2190 net657 net654 VDD VDD pmos w=2u l=1u
M2191 n2577 n2672 VDD VDD pmos w=2u l=1u
M2192 n2577 n2672 VSS VSS nmos w=1u l=1u
M2193 n2665 n2674 net658 VSS nmos w=1u l=1u
M2194 net658 n2673 VSS VSS nmos w=1u l=1u
M2195 n2665 n2674 VDD VDD pmos w=2u l=1u
M2196 n2665 n2673 VDD VDD pmos w=2u l=1u
M2197 net659 n2672 VSS VSS nmos w=1u l=1u
M2198 net660 n2576 VSS VSS nmos w=1u l=1u
M2199 n2674 net661 VSS VSS nmos w=1u l=1u
M2200 net661 n2672 net662 VSS nmos w=1u l=1u
M2201 net661 net659 net660 VSS nmos w=1u l=1u
M2202 net662 net660 VSS VSS nmos w=1u l=1u
M2203 net661 net659 net663 VDD pmos w=2u l=1u
M2204 net659 n2672 VDD VDD pmos w=2u l=1u
M2205 net660 n2672 net661 VDD pmos w=2u l=1u
M2206 net660 n2576 VDD VDD pmos w=2u l=1u
M2207 n2674 net661 VDD VDD pmos w=2u l=1u
M2208 net663 net660 VDD VDD pmos w=2u l=1u
M2209 n2672 N477 net664 VSS nmos w=1u l=1u
M2210 net664 N171 VSS VSS nmos w=1u l=1u
M2211 n2672 N477 VDD VDD pmos w=2u l=1u
M2212 n2672 N171 VDD VDD pmos w=2u l=1u
M2213 n2576 n2575 net665 VSS nmos w=1u l=1u
M2214 net665 n2675 VSS VSS nmos w=1u l=1u
M2215 n2576 n2575 VDD VDD pmos w=2u l=1u
M2216 n2576 n2675 VDD VDD pmos w=2u l=1u
M2217 n2575 n2677 net666 VSS nmos w=1u l=1u
M2218 net666 n2676 VSS VSS nmos w=1u l=1u
M2219 n2575 n2677 VDD VDD pmos w=2u l=1u
M2220 n2575 n2676 VDD VDD pmos w=2u l=1u
M2221 n2677 n2679 net667 VSS nmos w=1u l=1u
M2222 net667 n2678 VSS VSS nmos w=1u l=1u
M2223 n2677 n2679 VDD VDD pmos w=2u l=1u
M2224 n2677 n2678 VDD VDD pmos w=2u l=1u
M2225 n2678 net668 VSS VSS nmos w=1u l=1u
M2226 net668 n2680 VSS VSS nmos w=1u l=1u
M2227 net668 n2681 VSS VSS nmos w=1u l=1u
M2228 net668 n2681 net669 VDD pmos w=2u l=1u
M2229 n2678 net668 VDD VDD pmos w=2u l=1u
M2230 net669 n2680 VDD VDD pmos w=2u l=1u
M2231 net670 n2586 VSS VSS nmos w=1u l=1u
M2232 net671 n2587 VSS VSS nmos w=1u l=1u
M2233 n2676 net672 VSS VSS nmos w=1u l=1u
M2234 net672 n2586 net673 VSS nmos w=1u l=1u
M2235 net672 net670 net671 VSS nmos w=1u l=1u
M2236 net673 net671 VSS VSS nmos w=1u l=1u
M2237 net672 net670 net674 VDD pmos w=2u l=1u
M2238 net670 n2586 VDD VDD pmos w=2u l=1u
M2239 net671 n2586 net672 VDD pmos w=2u l=1u
M2240 net671 n2587 VDD VDD pmos w=2u l=1u
M2241 n2676 net672 VDD VDD pmos w=2u l=1u
M2242 net674 net671 VDD VDD pmos w=2u l=1u
M2243 n2587 n2682 VDD VDD pmos w=2u l=1u
M2244 n2587 n2682 VSS VSS nmos w=1u l=1u
M2245 n2675 n2684 net675 VSS nmos w=1u l=1u
M2246 net675 n2683 VSS VSS nmos w=1u l=1u
M2247 n2675 n2684 VDD VDD pmos w=2u l=1u
M2248 n2675 n2683 VDD VDD pmos w=2u l=1u
M2249 net676 n2682 VSS VSS nmos w=1u l=1u
M2250 net677 n2586 VSS VSS nmos w=1u l=1u
M2251 n2684 net678 VSS VSS nmos w=1u l=1u
M2252 net678 n2682 net679 VSS nmos w=1u l=1u
M2253 net678 net676 net677 VSS nmos w=1u l=1u
M2254 net679 net677 VSS VSS nmos w=1u l=1u
M2255 net678 net676 net680 VDD pmos w=2u l=1u
M2256 net676 n2682 VDD VDD pmos w=2u l=1u
M2257 net677 n2682 net678 VDD pmos w=2u l=1u
M2258 net677 n2586 VDD VDD pmos w=2u l=1u
M2259 n2684 net678 VDD VDD pmos w=2u l=1u
M2260 net680 net677 VDD VDD pmos w=2u l=1u
M2261 n2682 N460 net681 VSS nmos w=1u l=1u
M2262 net681 N188 VSS VSS nmos w=1u l=1u
M2263 n2682 N460 VDD VDD pmos w=2u l=1u
M2264 n2682 N188 VDD VDD pmos w=2u l=1u
M2265 n2586 n2585 net682 VSS nmos w=1u l=1u
M2266 net682 n2685 VSS VSS nmos w=1u l=1u
M2267 n2586 n2585 VDD VDD pmos w=2u l=1u
M2268 n2586 n2685 VDD VDD pmos w=2u l=1u
M2269 n2585 n2687 net683 VSS nmos w=1u l=1u
M2270 net683 n2686 VSS VSS nmos w=1u l=1u
M2271 n2585 n2687 VDD VDD pmos w=2u l=1u
M2272 n2585 n2686 VDD VDD pmos w=2u l=1u
M2273 n2687 n2689 net684 VSS nmos w=1u l=1u
M2274 net684 n2688 VSS VSS nmos w=1u l=1u
M2275 n2687 n2689 VDD VDD pmos w=2u l=1u
M2276 n2687 n2688 VDD VDD pmos w=2u l=1u
M2277 n2688 net685 VSS VSS nmos w=1u l=1u
M2278 net685 n2690 VSS VSS nmos w=1u l=1u
M2279 net685 n2691 VSS VSS nmos w=1u l=1u
M2280 net685 n2691 net686 VDD pmos w=2u l=1u
M2281 n2688 net685 VDD VDD pmos w=2u l=1u
M2282 net686 n2690 VDD VDD pmos w=2u l=1u
M2283 net687 n2596 VSS VSS nmos w=1u l=1u
M2284 net688 n2597 VSS VSS nmos w=1u l=1u
M2285 n2686 net689 VSS VSS nmos w=1u l=1u
M2286 net689 n2596 net690 VSS nmos w=1u l=1u
M2287 net689 net687 net688 VSS nmos w=1u l=1u
M2288 net690 net688 VSS VSS nmos w=1u l=1u
M2289 net689 net687 net691 VDD pmos w=2u l=1u
M2290 net687 n2596 VDD VDD pmos w=2u l=1u
M2291 net688 n2596 net689 VDD pmos w=2u l=1u
M2292 net688 n2597 VDD VDD pmos w=2u l=1u
M2293 n2686 net689 VDD VDD pmos w=2u l=1u
M2294 net691 net688 VDD VDD pmos w=2u l=1u
M2295 n2597 n2692 VDD VDD pmos w=2u l=1u
M2296 n2597 n2692 VSS VSS nmos w=1u l=1u
M2297 n2685 n2694 net692 VSS nmos w=1u l=1u
M2298 net692 n2693 VSS VSS nmos w=1u l=1u
M2299 n2685 n2694 VDD VDD pmos w=2u l=1u
M2300 n2685 n2693 VDD VDD pmos w=2u l=1u
M2301 net693 n2692 VSS VSS nmos w=1u l=1u
M2302 net694 n2596 VSS VSS nmos w=1u l=1u
M2303 n2694 net695 VSS VSS nmos w=1u l=1u
M2304 net695 n2692 net696 VSS nmos w=1u l=1u
M2305 net695 net693 net694 VSS nmos w=1u l=1u
M2306 net696 net694 VSS VSS nmos w=1u l=1u
M2307 net695 net693 net697 VDD pmos w=2u l=1u
M2308 net693 n2692 VDD VDD pmos w=2u l=1u
M2309 net694 n2692 net695 VDD pmos w=2u l=1u
M2310 net694 n2596 VDD VDD pmos w=2u l=1u
M2311 n2694 net695 VDD VDD pmos w=2u l=1u
M2312 net697 net694 VDD VDD pmos w=2u l=1u
M2313 n2692 N443 net698 VSS nmos w=1u l=1u
M2314 net698 N205 VSS VSS nmos w=1u l=1u
M2315 n2692 N443 VDD VDD pmos w=2u l=1u
M2316 n2692 N205 VDD VDD pmos w=2u l=1u
M2317 n2596 n2595 net699 VSS nmos w=1u l=1u
M2318 net699 n2695 VSS VSS nmos w=1u l=1u
M2319 n2596 n2595 VDD VDD pmos w=2u l=1u
M2320 n2596 n2695 VDD VDD pmos w=2u l=1u
M2321 n2595 n2697 net700 VSS nmos w=1u l=1u
M2322 net700 n2696 VSS VSS nmos w=1u l=1u
M2323 n2595 n2697 VDD VDD pmos w=2u l=1u
M2324 n2595 n2696 VDD VDD pmos w=2u l=1u
M2325 n2697 n2699 net701 VSS nmos w=1u l=1u
M2326 net701 n2698 VSS VSS nmos w=1u l=1u
M2327 n2697 n2699 VDD VDD pmos w=2u l=1u
M2328 n2697 n2698 VDD VDD pmos w=2u l=1u
M2329 n2698 n2701 net702 VSS nmos w=1u l=1u
M2330 net702 n2700 VSS VSS nmos w=1u l=1u
M2331 n2698 n2701 VDD VDD pmos w=2u l=1u
M2332 n2698 n2700 VDD VDD pmos w=2u l=1u
M2333 net703 n2607 VSS VSS nmos w=1u l=1u
M2334 net704 n2608 VSS VSS nmos w=1u l=1u
M2335 n2696 net705 VSS VSS nmos w=1u l=1u
M2336 net705 n2607 net706 VSS nmos w=1u l=1u
M2337 net705 net703 net704 VSS nmos w=1u l=1u
M2338 net706 net704 VSS VSS nmos w=1u l=1u
M2339 net705 net703 net707 VDD pmos w=2u l=1u
M2340 net703 n2607 VDD VDD pmos w=2u l=1u
M2341 net704 n2607 net705 VDD pmos w=2u l=1u
M2342 net704 n2608 VDD VDD pmos w=2u l=1u
M2343 n2696 net705 VDD VDD pmos w=2u l=1u
M2344 net707 net704 VDD VDD pmos w=2u l=1u
M2345 n2607 n2702 VDD VDD pmos w=2u l=1u
M2346 n2607 n2702 VSS VSS nmos w=1u l=1u
M2347 n2695 n2704 net708 VSS nmos w=1u l=1u
M2348 net708 n2703 VSS VSS nmos w=1u l=1u
M2349 n2695 n2704 VDD VDD pmos w=2u l=1u
M2350 n2695 n2703 VDD VDD pmos w=2u l=1u
M2351 net709 n2608 VSS VSS nmos w=1u l=1u
M2352 net710 n2702 VSS VSS nmos w=1u l=1u
M2353 n2704 net711 VSS VSS nmos w=1u l=1u
M2354 net711 n2608 net712 VSS nmos w=1u l=1u
M2355 net711 net709 net710 VSS nmos w=1u l=1u
M2356 net712 net710 VSS VSS nmos w=1u l=1u
M2357 net711 net709 net713 VDD pmos w=2u l=1u
M2358 net709 n2608 VDD VDD pmos w=2u l=1u
M2359 net710 n2608 net711 VDD pmos w=2u l=1u
M2360 net710 n2702 VDD VDD pmos w=2u l=1u
M2361 n2704 net711 VDD VDD pmos w=2u l=1u
M2362 net713 net710 VDD VDD pmos w=2u l=1u
M2363 n2608 N426 net714 VSS nmos w=1u l=1u
M2364 net714 N222 VSS VSS nmos w=1u l=1u
M2365 n2608 N426 VDD VDD pmos w=2u l=1u
M2366 n2608 N222 VDD VDD pmos w=2u l=1u
M2367 n2702 n2605 net715 VSS nmos w=1u l=1u
M2368 net715 n2705 VSS VSS nmos w=1u l=1u
M2369 n2702 n2605 VDD VDD pmos w=2u l=1u
M2370 n2702 n2705 VDD VDD pmos w=2u l=1u
M2371 n2605 n2707 net716 VSS nmos w=1u l=1u
M2372 net716 n2706 VSS VSS nmos w=1u l=1u
M2373 n2605 n2707 VDD VDD pmos w=2u l=1u
M2374 n2605 n2706 VDD VDD pmos w=2u l=1u
M2375 n2707 n2709 net717 VSS nmos w=1u l=1u
M2376 net717 n2708 VSS VSS nmos w=1u l=1u
M2377 n2707 n2709 VDD VDD pmos w=2u l=1u
M2378 n2707 n2708 VDD VDD pmos w=2u l=1u
M2379 n2705 n2708 net718 VSS nmos w=1u l=1u
M2380 net718 n2710 VSS VSS nmos w=1u l=1u
M2381 n2705 n2708 VDD VDD pmos w=2u l=1u
M2382 n2705 n2710 VDD VDD pmos w=2u l=1u
M2383 n2708 n2712 net719 VSS nmos w=1u l=1u
M2384 net719 n2711 VSS VSS nmos w=1u l=1u
M2385 n2708 n2712 VDD VDD pmos w=2u l=1u
M2386 n2708 n2711 VDD VDD pmos w=2u l=1u
M2387 n2710 n2706 VSS VSS nmos w=1u l=1u
M2388 n2710 n2713 VSS VSS nmos w=1u l=1u
M2389 n2710 n2706 net720 VDD pmos w=2u l=1u
M2390 net720 n2713 VDD VDD pmos w=2u l=1u
M2391 n2706 net721 VSS VSS nmos w=1u l=1u
M2392 net722 n2714 VSS VSS nmos w=1u l=1u
M2393 net721 n2620 net722 VSS nmos w=1u l=1u
M2394 net721 n2714 VDD VDD pmos w=2u l=1u
M2395 net721 n2620 VDD VDD pmos w=2u l=1u
M2396 n2706 net721 VDD VDD pmos w=2u l=1u
M2397 n2714 N409 net723 VSS nmos w=1u l=1u
M2398 net723 n2715 VSS VSS nmos w=1u l=1u
M2399 n2714 N409 VDD VDD pmos w=2u l=1u
M2400 n2714 n2715 VDD VDD pmos w=2u l=1u
M2401 n2715 n2717 VSS VSS nmos w=1u l=1u
M2402 n2715 n2716 VSS VSS nmos w=1u l=1u
M2403 n2715 n2717 net724 VDD pmos w=2u l=1u
M2404 net724 n2716 VDD VDD pmos w=2u l=1u
M2405 n2717 n2719 VSS VSS nmos w=1u l=1u
M2406 n2717 n2718 VSS VSS nmos w=1u l=1u
M2407 n2717 n2719 net725 VDD pmos w=2u l=1u
M2408 net725 n2718 VDD VDD pmos w=2u l=1u
M2409 n2719 n2270 net726 VSS nmos w=1u l=1u
M2410 net726 n2720 VSS VSS nmos w=1u l=1u
M2411 n2719 n2270 VDD VDD pmos w=2u l=1u
M2412 n2719 n2720 VDD VDD pmos w=2u l=1u
M2413 n2720 n2721 net727 VSS nmos w=1u l=1u
M2414 net727 N239 VSS VSS nmos w=1u l=1u
M2415 n2720 n2721 VDD VDD pmos w=2u l=1u
M2416 n2720 N239 VDD VDD pmos w=2u l=1u
M2417 n2718 n2623 VDD VDD pmos w=2u l=1u
M2418 n2718 n2623 VSS VSS nmos w=1u l=1u
M2419 n2716 n2623 VSS VSS nmos w=1u l=1u
M2420 n2716 N392 VSS VSS nmos w=1u l=1u
M2421 n2716 n2623 net728 VDD pmos w=2u l=1u
M2422 net728 N392 VDD VDD pmos w=2u l=1u
M2423 n2620 n2723 net729 VSS nmos w=1u l=1u
M2424 net729 n2722 VSS VSS nmos w=1u l=1u
M2425 n2620 n2723 VDD VDD pmos w=2u l=1u
M2426 n2620 n2722 VDD VDD pmos w=2u l=1u
M2427 n2723 N239 net730 VSS nmos w=1u l=1u
M2428 net730 N409 VSS VSS nmos w=1u l=1u
M2429 n2723 N239 VDD VDD pmos w=2u l=1u
M2430 n2723 N409 VDD VDD pmos w=2u l=1u
M2431 net731 n2622 VSS VSS nmos w=1u l=1u
M2432 net732 n2623 VSS VSS nmos w=1u l=1u
M2433 n2722 net733 VSS VSS nmos w=1u l=1u
M2434 net733 n2622 net734 VSS nmos w=1u l=1u
M2435 net733 net731 net732 VSS nmos w=1u l=1u
M2436 net734 net732 VSS VSS nmos w=1u l=1u
M2437 net733 net731 net735 VDD pmos w=2u l=1u
M2438 net731 n2622 VDD VDD pmos w=2u l=1u
M2439 net732 n2622 net733 VDD pmos w=2u l=1u
M2440 net732 n2623 VDD VDD pmos w=2u l=1u
M2441 n2722 net733 VDD VDD pmos w=2u l=1u
M2442 net735 net732 VDD VDD pmos w=2u l=1u
M2443 n2622 N256 net736 VSS nmos w=1u l=1u
M2444 net736 N392 VSS VSS nmos w=1u l=1u
M2445 n2622 N256 VDD VDD pmos w=2u l=1u
M2446 n2622 N392 VDD VDD pmos w=2u l=1u
M2447 n2623 n2725 net737 VSS nmos w=1u l=1u
M2448 net737 n2724 VSS VSS nmos w=1u l=1u
M2449 n2623 n2725 VDD VDD pmos w=2u l=1u
M2450 n2623 n2724 VDD VDD pmos w=2u l=1u
M2451 n2725 n2727 net738 VSS nmos w=1u l=1u
M2452 net738 n2726 VSS VSS nmos w=1u l=1u
M2453 n2725 n2727 VDD VDD pmos w=2u l=1u
M2454 n2725 n2726 VDD VDD pmos w=2u l=1u
M2455 n2713 n2709 VDD VDD pmos w=2u l=1u
M2456 n2713 n2709 VSS VSS nmos w=1u l=1u
M2457 n2703 n2729 VSS VSS nmos w=1u l=1u
M2458 n2703 n2728 VSS VSS nmos w=1u l=1u
M2459 n2703 n2729 net739 VDD pmos w=2u l=1u
M2460 net739 n2728 VDD VDD pmos w=2u l=1u
M2461 n2729 net740 VSS VSS nmos w=1u l=1u
M2462 net741 n2700 VSS VSS nmos w=1u l=1u
M2463 net740 n2701 net741 VSS nmos w=1u l=1u
M2464 net740 n2700 VDD VDD pmos w=2u l=1u
M2465 net740 n2701 VDD VDD pmos w=2u l=1u
M2466 n2729 net740 VDD VDD pmos w=2u l=1u
M2467 n2728 n2699 VDD VDD pmos w=2u l=1u
M2468 n2728 n2699 VSS VSS nmos w=1u l=1u
M2469 n2693 n2731 VSS VSS nmos w=1u l=1u
M2470 n2693 n2730 VSS VSS nmos w=1u l=1u
M2471 n2693 n2731 net742 VDD pmos w=2u l=1u
M2472 net742 n2730 VDD VDD pmos w=2u l=1u
M2473 n2731 n2690 VSS VSS nmos w=1u l=1u
M2474 n2731 n2691 VSS VSS nmos w=1u l=1u
M2475 n2731 n2690 net743 VDD pmos w=2u l=1u
M2476 net743 n2691 VDD VDD pmos w=2u l=1u
M2477 n2730 n2689 VDD VDD pmos w=2u l=1u
M2478 n2730 n2689 VSS VSS nmos w=1u l=1u
M2479 n2683 n2733 VSS VSS nmos w=1u l=1u
M2480 n2683 n2732 VSS VSS nmos w=1u l=1u
M2481 n2683 n2733 net744 VDD pmos w=2u l=1u
M2482 net744 n2732 VDD VDD pmos w=2u l=1u
M2483 n2733 n2680 VSS VSS nmos w=1u l=1u
M2484 n2733 n2681 VSS VSS nmos w=1u l=1u
M2485 n2733 n2680 net745 VDD pmos w=2u l=1u
M2486 net745 n2681 VDD VDD pmos w=2u l=1u
M2487 n2732 n2679 VDD VDD pmos w=2u l=1u
M2488 n2732 n2679 VSS VSS nmos w=1u l=1u
M2489 n2673 n2735 VSS VSS nmos w=1u l=1u
M2490 n2673 n2734 VSS VSS nmos w=1u l=1u
M2491 n2673 n2735 net746 VDD pmos w=2u l=1u
M2492 net746 n2734 VDD VDD pmos w=2u l=1u
M2493 n2735 n2670 VSS VSS nmos w=1u l=1u
M2494 n2735 n2671 VSS VSS nmos w=1u l=1u
M2495 n2735 n2670 net747 VDD pmos w=2u l=1u
M2496 net747 n2671 VDD VDD pmos w=2u l=1u
M2497 n2734 n2669 VDD VDD pmos w=2u l=1u
M2498 n2734 n2669 VSS VSS nmos w=1u l=1u
M2499 n2663 n2737 VSS VSS nmos w=1u l=1u
M2500 n2663 n2736 VSS VSS nmos w=1u l=1u
M2501 n2663 n2737 net748 VDD pmos w=2u l=1u
M2502 net748 n2736 VDD VDD pmos w=2u l=1u
M2503 n2737 n2660 VSS VSS nmos w=1u l=1u
M2504 n2737 n2661 VSS VSS nmos w=1u l=1u
M2505 n2737 n2660 net749 VDD pmos w=2u l=1u
M2506 net749 n2661 VDD VDD pmos w=2u l=1u
M2507 n2736 n2659 VDD VDD pmos w=2u l=1u
M2508 n2736 n2659 VSS VSS nmos w=1u l=1u
M2509 n2653 n2739 VSS VSS nmos w=1u l=1u
M2510 n2653 n2738 VSS VSS nmos w=1u l=1u
M2511 n2653 n2739 net750 VDD pmos w=2u l=1u
M2512 net750 n2738 VDD VDD pmos w=2u l=1u
M2513 n2739 n2650 VSS VSS nmos w=1u l=1u
M2514 n2739 n2651 VSS VSS nmos w=1u l=1u
M2515 n2739 n2650 net751 VDD pmos w=2u l=1u
M2516 net751 n2651 VDD VDD pmos w=2u l=1u
M2517 n2738 n2649 VDD VDD pmos w=2u l=1u
M2518 n2738 n2649 VSS VSS nmos w=1u l=1u
M2519 n2550 N528 net752 VSS nmos w=1u l=1u
M2520 net752 N120 VSS VSS nmos w=1u l=1u
M2521 n2550 N528 VDD VDD pmos w=2u l=1u
M2522 n2550 N120 VDD VDD pmos w=2u l=1u
M2523 N6200 n2740 net753 VSS nmos w=1u l=1u
M2524 net753 n2638 VSS VSS nmos w=1u l=1u
M2525 N6200 n2740 VDD VDD pmos w=2u l=1u
M2526 N6200 n2638 VDD VDD pmos w=2u l=1u
M2527 n2740 net754 VSS VSS nmos w=1u l=1u
M2528 net754 n2741 VSS VSS nmos w=1u l=1u
M2529 net754 n2742 VSS VSS nmos w=1u l=1u
M2530 net754 n2742 net755 VDD pmos w=2u l=1u
M2531 n2740 net754 VDD VDD pmos w=2u l=1u
M2532 net755 n2741 VDD VDD pmos w=2u l=1u
M2533 n2638 n2742 net756 VSS nmos w=1u l=1u
M2534 net756 n2741 VSS VSS nmos w=1u l=1u
M2535 n2638 n2742 VDD VDD pmos w=2u l=1u
M2536 n2638 n2741 VDD VDD pmos w=2u l=1u
M2537 n2742 n2744 net757 VSS nmos w=1u l=1u
M2538 net757 n2743 VSS VSS nmos w=1u l=1u
M2539 n2742 n2744 VDD VDD pmos w=2u l=1u
M2540 n2742 n2743 VDD VDD pmos w=2u l=1u
M2541 n2743 n2746 net758 VSS nmos w=1u l=1u
M2542 net758 n2745 VSS VSS nmos w=1u l=1u
M2543 n2743 n2746 VDD VDD pmos w=2u l=1u
M2544 n2743 n2745 VDD VDD pmos w=2u l=1u
M2545 net759 n2640 VSS VSS nmos w=1u l=1u
M2546 net760 n2639 VSS VSS nmos w=1u l=1u
M2547 n2741 net761 VSS VSS nmos w=1u l=1u
M2548 net761 n2640 net762 VSS nmos w=1u l=1u
M2549 net761 net759 net760 VSS nmos w=1u l=1u
M2550 net762 net760 VSS VSS nmos w=1u l=1u
M2551 net761 net759 net763 VDD pmos w=2u l=1u
M2552 net759 n2640 VDD VDD pmos w=2u l=1u
M2553 net760 n2640 net761 VDD pmos w=2u l=1u
M2554 net760 n2639 VDD VDD pmos w=2u l=1u
M2555 n2741 net761 VDD VDD pmos w=2u l=1u
M2556 net763 net760 VDD VDD pmos w=2u l=1u
M2557 n2640 n2748 net764 VSS nmos w=1u l=1u
M2558 net764 n2747 VSS VSS nmos w=1u l=1u
M2559 n2640 n2748 VDD VDD pmos w=2u l=1u
M2560 n2640 n2747 VDD VDD pmos w=2u l=1u
M2561 n2747 n2750 net765 VSS nmos w=1u l=1u
M2562 net765 n2749 VSS VSS nmos w=1u l=1u
M2563 n2747 n2750 VDD VDD pmos w=2u l=1u
M2564 n2747 n2749 VDD VDD pmos w=2u l=1u
M2565 net766 n2643 VSS VSS nmos w=1u l=1u
M2566 net767 n2644 VSS VSS nmos w=1u l=1u
M2567 n2639 net768 VSS VSS nmos w=1u l=1u
M2568 net768 n2643 net769 VSS nmos w=1u l=1u
M2569 net768 net766 net767 VSS nmos w=1u l=1u
M2570 net769 net767 VSS VSS nmos w=1u l=1u
M2571 net768 net766 net770 VDD pmos w=2u l=1u
M2572 net766 n2643 VDD VDD pmos w=2u l=1u
M2573 net767 n2643 net768 VDD pmos w=2u l=1u
M2574 net767 n2644 VDD VDD pmos w=2u l=1u
M2575 n2639 net768 VDD VDD pmos w=2u l=1u
M2576 net770 net767 VDD VDD pmos w=2u l=1u
M2577 n2643 net771 VSS VSS nmos w=1u l=1u
M2578 net772 n2642 VSS VSS nmos w=1u l=1u
M2579 net771 n2751 net772 VSS nmos w=1u l=1u
M2580 net771 n2642 VDD VDD pmos w=2u l=1u
M2581 net771 n2751 VDD VDD pmos w=2u l=1u
M2582 n2643 net771 VDD VDD pmos w=2u l=1u
M2583 n2642 n2753 net773 VSS nmos w=1u l=1u
M2584 net773 n2752 VSS VSS nmos w=1u l=1u
M2585 n2642 n2753 VDD VDD pmos w=2u l=1u
M2586 n2642 n2752 VDD VDD pmos w=2u l=1u
M2587 n2753 n2755 net774 VSS nmos w=1u l=1u
M2588 net774 n2754 VSS VSS nmos w=1u l=1u
M2589 n2753 n2755 VDD VDD pmos w=2u l=1u
M2590 n2753 n2754 VDD VDD pmos w=2u l=1u
M2591 n2754 net775 VSS VSS nmos w=1u l=1u
M2592 net775 n2756 VSS VSS nmos w=1u l=1u
M2593 net775 n2757 VSS VSS nmos w=1u l=1u
M2594 net775 n2757 net776 VDD pmos w=2u l=1u
M2595 n2754 net775 VDD VDD pmos w=2u l=1u
M2596 net776 n2756 VDD VDD pmos w=2u l=1u
M2597 net777 n2650 VSS VSS nmos w=1u l=1u
M2598 net778 n2651 VSS VSS nmos w=1u l=1u
M2599 n2752 net779 VSS VSS nmos w=1u l=1u
M2600 net779 n2650 net780 VSS nmos w=1u l=1u
M2601 net779 net777 net778 VSS nmos w=1u l=1u
M2602 net780 net778 VSS VSS nmos w=1u l=1u
M2603 net779 net777 net781 VDD pmos w=2u l=1u
M2604 net777 n2650 VDD VDD pmos w=2u l=1u
M2605 net778 n2650 net779 VDD pmos w=2u l=1u
M2606 net778 n2651 VDD VDD pmos w=2u l=1u
M2607 n2752 net779 VDD VDD pmos w=2u l=1u
M2608 net781 net778 VDD VDD pmos w=2u l=1u
M2609 n2651 n2758 VDD VDD pmos w=2u l=1u
M2610 n2651 n2758 VSS VSS nmos w=1u l=1u
M2611 n2751 n2760 net782 VSS nmos w=1u l=1u
M2612 net782 n2759 VSS VSS nmos w=1u l=1u
M2613 n2751 n2760 VDD VDD pmos w=2u l=1u
M2614 n2751 n2759 VDD VDD pmos w=2u l=1u
M2615 net783 n2758 VSS VSS nmos w=1u l=1u
M2616 net784 n2650 VSS VSS nmos w=1u l=1u
M2617 n2760 net785 VSS VSS nmos w=1u l=1u
M2618 net785 n2758 net786 VSS nmos w=1u l=1u
M2619 net785 net783 net784 VSS nmos w=1u l=1u
M2620 net786 net784 VSS VSS nmos w=1u l=1u
M2621 net785 net783 net787 VDD pmos w=2u l=1u
M2622 net783 n2758 VDD VDD pmos w=2u l=1u
M2623 net784 n2758 net785 VDD pmos w=2u l=1u
M2624 net784 n2650 VDD VDD pmos w=2u l=1u
M2625 n2760 net785 VDD VDD pmos w=2u l=1u
M2626 net787 net784 VDD VDD pmos w=2u l=1u
M2627 n2758 N511 net788 VSS nmos w=1u l=1u
M2628 net788 N120 VSS VSS nmos w=1u l=1u
M2629 n2758 N511 VDD VDD pmos w=2u l=1u
M2630 n2758 N120 VDD VDD pmos w=2u l=1u
M2631 n2650 n2649 net789 VSS nmos w=1u l=1u
M2632 net789 n2761 VSS VSS nmos w=1u l=1u
M2633 n2650 n2649 VDD VDD pmos w=2u l=1u
M2634 n2650 n2761 VDD VDD pmos w=2u l=1u
M2635 n2649 n2763 net790 VSS nmos w=1u l=1u
M2636 net790 n2762 VSS VSS nmos w=1u l=1u
M2637 n2649 n2763 VDD VDD pmos w=2u l=1u
M2638 n2649 n2762 VDD VDD pmos w=2u l=1u
M2639 n2763 n2765 net791 VSS nmos w=1u l=1u
M2640 net791 n2764 VSS VSS nmos w=1u l=1u
M2641 n2763 n2765 VDD VDD pmos w=2u l=1u
M2642 n2763 n2764 VDD VDD pmos w=2u l=1u
M2643 n2764 net792 VSS VSS nmos w=1u l=1u
M2644 net792 n2766 VSS VSS nmos w=1u l=1u
M2645 net792 n2767 VSS VSS nmos w=1u l=1u
M2646 net792 n2767 net793 VDD pmos w=2u l=1u
M2647 n2764 net792 VDD VDD pmos w=2u l=1u
M2648 net793 n2766 VDD VDD pmos w=2u l=1u
M2649 net794 n2660 VSS VSS nmos w=1u l=1u
M2650 net795 n2661 VSS VSS nmos w=1u l=1u
M2651 n2762 net796 VSS VSS nmos w=1u l=1u
M2652 net796 n2660 net797 VSS nmos w=1u l=1u
M2653 net796 net794 net795 VSS nmos w=1u l=1u
M2654 net797 net795 VSS VSS nmos w=1u l=1u
M2655 net796 net794 net798 VDD pmos w=2u l=1u
M2656 net794 n2660 VDD VDD pmos w=2u l=1u
M2657 net795 n2660 net796 VDD pmos w=2u l=1u
M2658 net795 n2661 VDD VDD pmos w=2u l=1u
M2659 n2762 net796 VDD VDD pmos w=2u l=1u
M2660 net798 net795 VDD VDD pmos w=2u l=1u
M2661 n2661 n2768 VDD VDD pmos w=2u l=1u
M2662 n2661 n2768 VSS VSS nmos w=1u l=1u
M2663 n2761 n2770 net799 VSS nmos w=1u l=1u
M2664 net799 n2769 VSS VSS nmos w=1u l=1u
M2665 n2761 n2770 VDD VDD pmos w=2u l=1u
M2666 n2761 n2769 VDD VDD pmos w=2u l=1u
M2667 net800 n2768 VSS VSS nmos w=1u l=1u
M2668 net801 n2660 VSS VSS nmos w=1u l=1u
M2669 n2770 net802 VSS VSS nmos w=1u l=1u
M2670 net802 n2768 net803 VSS nmos w=1u l=1u
M2671 net802 net800 net801 VSS nmos w=1u l=1u
M2672 net803 net801 VSS VSS nmos w=1u l=1u
M2673 net802 net800 net804 VDD pmos w=2u l=1u
M2674 net800 n2768 VDD VDD pmos w=2u l=1u
M2675 net801 n2768 net802 VDD pmos w=2u l=1u
M2676 net801 n2660 VDD VDD pmos w=2u l=1u
M2677 n2770 net802 VDD VDD pmos w=2u l=1u
M2678 net804 net801 VDD VDD pmos w=2u l=1u
M2679 n2768 N494 net805 VSS nmos w=1u l=1u
M2680 net805 N137 VSS VSS nmos w=1u l=1u
M2681 n2768 N494 VDD VDD pmos w=2u l=1u
M2682 n2768 N137 VDD VDD pmos w=2u l=1u
M2683 n2660 n2659 net806 VSS nmos w=1u l=1u
M2684 net806 n2771 VSS VSS nmos w=1u l=1u
M2685 n2660 n2659 VDD VDD pmos w=2u l=1u
M2686 n2660 n2771 VDD VDD pmos w=2u l=1u
M2687 n2659 n2773 net807 VSS nmos w=1u l=1u
M2688 net807 n2772 VSS VSS nmos w=1u l=1u
M2689 n2659 n2773 VDD VDD pmos w=2u l=1u
M2690 n2659 n2772 VDD VDD pmos w=2u l=1u
M2691 n2773 n2775 net808 VSS nmos w=1u l=1u
M2692 net808 n2774 VSS VSS nmos w=1u l=1u
M2693 n2773 n2775 VDD VDD pmos w=2u l=1u
M2694 n2773 n2774 VDD VDD pmos w=2u l=1u
M2695 n2774 net809 VSS VSS nmos w=1u l=1u
M2696 net809 n2776 VSS VSS nmos w=1u l=1u
M2697 net809 n2777 VSS VSS nmos w=1u l=1u
M2698 net809 n2777 net810 VDD pmos w=2u l=1u
M2699 n2774 net809 VDD VDD pmos w=2u l=1u
M2700 net810 n2776 VDD VDD pmos w=2u l=1u
M2701 net811 n2670 VSS VSS nmos w=1u l=1u
M2702 net812 n2671 VSS VSS nmos w=1u l=1u
M2703 n2772 net813 VSS VSS nmos w=1u l=1u
M2704 net813 n2670 net814 VSS nmos w=1u l=1u
M2705 net813 net811 net812 VSS nmos w=1u l=1u
M2706 net814 net812 VSS VSS nmos w=1u l=1u
M2707 net813 net811 net815 VDD pmos w=2u l=1u
M2708 net811 n2670 VDD VDD pmos w=2u l=1u
M2709 net812 n2670 net813 VDD pmos w=2u l=1u
M2710 net812 n2671 VDD VDD pmos w=2u l=1u
M2711 n2772 net813 VDD VDD pmos w=2u l=1u
M2712 net815 net812 VDD VDD pmos w=2u l=1u
M2713 n2671 n2778 VDD VDD pmos w=2u l=1u
M2714 n2671 n2778 VSS VSS nmos w=1u l=1u
M2715 n2771 n2780 net816 VSS nmos w=1u l=1u
M2716 net816 n2779 VSS VSS nmos w=1u l=1u
M2717 n2771 n2780 VDD VDD pmos w=2u l=1u
M2718 n2771 n2779 VDD VDD pmos w=2u l=1u
M2719 net817 n2778 VSS VSS nmos w=1u l=1u
M2720 net818 n2670 VSS VSS nmos w=1u l=1u
M2721 n2780 net819 VSS VSS nmos w=1u l=1u
M2722 net819 n2778 net820 VSS nmos w=1u l=1u
M2723 net819 net817 net818 VSS nmos w=1u l=1u
M2724 net820 net818 VSS VSS nmos w=1u l=1u
M2725 net819 net817 net821 VDD pmos w=2u l=1u
M2726 net817 n2778 VDD VDD pmos w=2u l=1u
M2727 net818 n2778 net819 VDD pmos w=2u l=1u
M2728 net818 n2670 VDD VDD pmos w=2u l=1u
M2729 n2780 net819 VDD VDD pmos w=2u l=1u
M2730 net821 net818 VDD VDD pmos w=2u l=1u
M2731 n2778 N477 net822 VSS nmos w=1u l=1u
M2732 net822 N154 VSS VSS nmos w=1u l=1u
M2733 n2778 N477 VDD VDD pmos w=2u l=1u
M2734 n2778 N154 VDD VDD pmos w=2u l=1u
M2735 n2670 n2669 net823 VSS nmos w=1u l=1u
M2736 net823 n2781 VSS VSS nmos w=1u l=1u
M2737 n2670 n2669 VDD VDD pmos w=2u l=1u
M2738 n2670 n2781 VDD VDD pmos w=2u l=1u
M2739 n2669 n2783 net824 VSS nmos w=1u l=1u
M2740 net824 n2782 VSS VSS nmos w=1u l=1u
M2741 n2669 n2783 VDD VDD pmos w=2u l=1u
M2742 n2669 n2782 VDD VDD pmos w=2u l=1u
M2743 n2783 n2785 net825 VSS nmos w=1u l=1u
M2744 net825 n2784 VSS VSS nmos w=1u l=1u
M2745 n2783 n2785 VDD VDD pmos w=2u l=1u
M2746 n2783 n2784 VDD VDD pmos w=2u l=1u
M2747 n2784 net826 VSS VSS nmos w=1u l=1u
M2748 net826 n2786 VSS VSS nmos w=1u l=1u
M2749 net826 n2787 VSS VSS nmos w=1u l=1u
M2750 net826 n2787 net827 VDD pmos w=2u l=1u
M2751 n2784 net826 VDD VDD pmos w=2u l=1u
M2752 net827 n2786 VDD VDD pmos w=2u l=1u
M2753 net828 n2680 VSS VSS nmos w=1u l=1u
M2754 net829 n2681 VSS VSS nmos w=1u l=1u
M2755 n2782 net830 VSS VSS nmos w=1u l=1u
M2756 net830 n2680 net831 VSS nmos w=1u l=1u
M2757 net830 net828 net829 VSS nmos w=1u l=1u
M2758 net831 net829 VSS VSS nmos w=1u l=1u
M2759 net830 net828 net832 VDD pmos w=2u l=1u
M2760 net828 n2680 VDD VDD pmos w=2u l=1u
M2761 net829 n2680 net830 VDD pmos w=2u l=1u
M2762 net829 n2681 VDD VDD pmos w=2u l=1u
M2763 n2782 net830 VDD VDD pmos w=2u l=1u
M2764 net832 net829 VDD VDD pmos w=2u l=1u
M2765 n2681 n2788 VDD VDD pmos w=2u l=1u
M2766 n2681 n2788 VSS VSS nmos w=1u l=1u
M2767 n2781 n2790 net833 VSS nmos w=1u l=1u
M2768 net833 n2789 VSS VSS nmos w=1u l=1u
M2769 n2781 n2790 VDD VDD pmos w=2u l=1u
M2770 n2781 n2789 VDD VDD pmos w=2u l=1u
M2771 net834 n2788 VSS VSS nmos w=1u l=1u
M2772 net835 n2680 VSS VSS nmos w=1u l=1u
M2773 n2790 net836 VSS VSS nmos w=1u l=1u
M2774 net836 n2788 net837 VSS nmos w=1u l=1u
M2775 net836 net834 net835 VSS nmos w=1u l=1u
M2776 net837 net835 VSS VSS nmos w=1u l=1u
M2777 net836 net834 net838 VDD pmos w=2u l=1u
M2778 net834 n2788 VDD VDD pmos w=2u l=1u
M2779 net835 n2788 net836 VDD pmos w=2u l=1u
M2780 net835 n2680 VDD VDD pmos w=2u l=1u
M2781 n2790 net836 VDD VDD pmos w=2u l=1u
M2782 net838 net835 VDD VDD pmos w=2u l=1u
M2783 n2788 N460 net839 VSS nmos w=1u l=1u
M2784 net839 N171 VSS VSS nmos w=1u l=1u
M2785 n2788 N460 VDD VDD pmos w=2u l=1u
M2786 n2788 N171 VDD VDD pmos w=2u l=1u
M2787 n2680 n2679 net840 VSS nmos w=1u l=1u
M2788 net840 n2791 VSS VSS nmos w=1u l=1u
M2789 n2680 n2679 VDD VDD pmos w=2u l=1u
M2790 n2680 n2791 VDD VDD pmos w=2u l=1u
M2791 n2679 n2793 net841 VSS nmos w=1u l=1u
M2792 net841 n2792 VSS VSS nmos w=1u l=1u
M2793 n2679 n2793 VDD VDD pmos w=2u l=1u
M2794 n2679 n2792 VDD VDD pmos w=2u l=1u
M2795 n2793 n2795 net842 VSS nmos w=1u l=1u
M2796 net842 n2794 VSS VSS nmos w=1u l=1u
M2797 n2793 n2795 VDD VDD pmos w=2u l=1u
M2798 n2793 n2794 VDD VDD pmos w=2u l=1u
M2799 n2794 net843 VSS VSS nmos w=1u l=1u
M2800 net843 n2796 VSS VSS nmos w=1u l=1u
M2801 net843 n2797 VSS VSS nmos w=1u l=1u
M2802 net843 n2797 net844 VDD pmos w=2u l=1u
M2803 n2794 net843 VDD VDD pmos w=2u l=1u
M2804 net844 n2796 VDD VDD pmos w=2u l=1u
M2805 net845 n2690 VSS VSS nmos w=1u l=1u
M2806 net846 n2691 VSS VSS nmos w=1u l=1u
M2807 n2792 net847 VSS VSS nmos w=1u l=1u
M2808 net847 n2690 net848 VSS nmos w=1u l=1u
M2809 net847 net845 net846 VSS nmos w=1u l=1u
M2810 net848 net846 VSS VSS nmos w=1u l=1u
M2811 net847 net845 net849 VDD pmos w=2u l=1u
M2812 net845 n2690 VDD VDD pmos w=2u l=1u
M2813 net846 n2690 net847 VDD pmos w=2u l=1u
M2814 net846 n2691 VDD VDD pmos w=2u l=1u
M2815 n2792 net847 VDD VDD pmos w=2u l=1u
M2816 net849 net846 VDD VDD pmos w=2u l=1u
M2817 n2691 n2798 VDD VDD pmos w=2u l=1u
M2818 n2691 n2798 VSS VSS nmos w=1u l=1u
M2819 n2791 n2800 net850 VSS nmos w=1u l=1u
M2820 net850 n2799 VSS VSS nmos w=1u l=1u
M2821 n2791 n2800 VDD VDD pmos w=2u l=1u
M2822 n2791 n2799 VDD VDD pmos w=2u l=1u
M2823 net851 n2798 VSS VSS nmos w=1u l=1u
M2824 net852 n2690 VSS VSS nmos w=1u l=1u
M2825 n2800 net853 VSS VSS nmos w=1u l=1u
M2826 net853 n2798 net854 VSS nmos w=1u l=1u
M2827 net853 net851 net852 VSS nmos w=1u l=1u
M2828 net854 net852 VSS VSS nmos w=1u l=1u
M2829 net853 net851 net855 VDD pmos w=2u l=1u
M2830 net851 n2798 VDD VDD pmos w=2u l=1u
M2831 net852 n2798 net853 VDD pmos w=2u l=1u
M2832 net852 n2690 VDD VDD pmos w=2u l=1u
M2833 n2800 net853 VDD VDD pmos w=2u l=1u
M2834 net855 net852 VDD VDD pmos w=2u l=1u
M2835 n2798 N443 net856 VSS nmos w=1u l=1u
M2836 net856 N188 VSS VSS nmos w=1u l=1u
M2837 n2798 N443 VDD VDD pmos w=2u l=1u
M2838 n2798 N188 VDD VDD pmos w=2u l=1u
M2839 n2690 n2689 net857 VSS nmos w=1u l=1u
M2840 net857 n2801 VSS VSS nmos w=1u l=1u
M2841 n2690 n2689 VDD VDD pmos w=2u l=1u
M2842 n2690 n2801 VDD VDD pmos w=2u l=1u
M2843 n2689 n2803 net858 VSS nmos w=1u l=1u
M2844 net858 n2802 VSS VSS nmos w=1u l=1u
M2845 n2689 n2803 VDD VDD pmos w=2u l=1u
M2846 n2689 n2802 VDD VDD pmos w=2u l=1u
M2847 n2803 n2805 net859 VSS nmos w=1u l=1u
M2848 net859 n2804 VSS VSS nmos w=1u l=1u
M2849 n2803 n2805 VDD VDD pmos w=2u l=1u
M2850 n2803 n2804 VDD VDD pmos w=2u l=1u
M2851 n2804 net860 VSS VSS nmos w=1u l=1u
M2852 net860 n2806 VSS VSS nmos w=1u l=1u
M2853 net860 n2807 VSS VSS nmos w=1u l=1u
M2854 net860 n2807 net861 VDD pmos w=2u l=1u
M2855 n2804 net860 VDD VDD pmos w=2u l=1u
M2856 net861 n2806 VDD VDD pmos w=2u l=1u
M2857 net862 n2700 VSS VSS nmos w=1u l=1u
M2858 net863 n2701 VSS VSS nmos w=1u l=1u
M2859 n2802 net864 VSS VSS nmos w=1u l=1u
M2860 net864 n2700 net865 VSS nmos w=1u l=1u
M2861 net864 net862 net863 VSS nmos w=1u l=1u
M2862 net865 net863 VSS VSS nmos w=1u l=1u
M2863 net864 net862 net866 VDD pmos w=2u l=1u
M2864 net862 n2700 VDD VDD pmos w=2u l=1u
M2865 net863 n2700 net864 VDD pmos w=2u l=1u
M2866 net863 n2701 VDD VDD pmos w=2u l=1u
M2867 n2802 net864 VDD VDD pmos w=2u l=1u
M2868 net866 net863 VDD VDD pmos w=2u l=1u
M2869 n2700 n2808 VDD VDD pmos w=2u l=1u
M2870 n2700 n2808 VSS VSS nmos w=1u l=1u
M2871 n2801 n2810 net867 VSS nmos w=1u l=1u
M2872 net867 n2809 VSS VSS nmos w=1u l=1u
M2873 n2801 n2810 VDD VDD pmos w=2u l=1u
M2874 n2801 n2809 VDD VDD pmos w=2u l=1u
M2875 net868 n2701 VSS VSS nmos w=1u l=1u
M2876 net869 n2808 VSS VSS nmos w=1u l=1u
M2877 n2810 net870 VSS VSS nmos w=1u l=1u
M2878 net870 n2701 net871 VSS nmos w=1u l=1u
M2879 net870 net868 net869 VSS nmos w=1u l=1u
M2880 net871 net869 VSS VSS nmos w=1u l=1u
M2881 net870 net868 net872 VDD pmos w=2u l=1u
M2882 net868 n2701 VDD VDD pmos w=2u l=1u
M2883 net869 n2701 net870 VDD pmos w=2u l=1u
M2884 net869 n2808 VDD VDD pmos w=2u l=1u
M2885 n2810 net870 VDD VDD pmos w=2u l=1u
M2886 net872 net869 VDD VDD pmos w=2u l=1u
M2887 n2701 N426 net873 VSS nmos w=1u l=1u
M2888 net873 N205 VSS VSS nmos w=1u l=1u
M2889 n2701 N426 VDD VDD pmos w=2u l=1u
M2890 n2701 N205 VDD VDD pmos w=2u l=1u
M2891 n2808 n2699 net874 VSS nmos w=1u l=1u
M2892 net874 n2811 VSS VSS nmos w=1u l=1u
M2893 n2808 n2699 VDD VDD pmos w=2u l=1u
M2894 n2808 n2811 VDD VDD pmos w=2u l=1u
M2895 n2699 n2813 net875 VSS nmos w=1u l=1u
M2896 net875 n2812 VSS VSS nmos w=1u l=1u
M2897 n2699 n2813 VDD VDD pmos w=2u l=1u
M2898 n2699 n2812 VDD VDD pmos w=2u l=1u
M2899 n2813 n2815 net876 VSS nmos w=1u l=1u
M2900 net876 n2814 VSS VSS nmos w=1u l=1u
M2901 n2813 n2815 VDD VDD pmos w=2u l=1u
M2902 n2813 n2814 VDD VDD pmos w=2u l=1u
M2903 n2814 net877 VSS VSS nmos w=1u l=1u
M2904 net877 n2816 VSS VSS nmos w=1u l=1u
M2905 net877 n2817 VSS VSS nmos w=1u l=1u
M2906 net877 n2817 net878 VDD pmos w=2u l=1u
M2907 n2814 net877 VDD VDD pmos w=2u l=1u
M2908 net878 n2816 VDD VDD pmos w=2u l=1u
M2909 net879 n2711 VSS VSS nmos w=1u l=1u
M2910 net880 n2712 VSS VSS nmos w=1u l=1u
M2911 n2812 net881 VSS VSS nmos w=1u l=1u
M2912 net881 n2711 net882 VSS nmos w=1u l=1u
M2913 net881 net879 net880 VSS nmos w=1u l=1u
M2914 net882 net880 VSS VSS nmos w=1u l=1u
M2915 net881 net879 net883 VDD pmos w=2u l=1u
M2916 net879 n2711 VDD VDD pmos w=2u l=1u
M2917 net880 n2711 net881 VDD pmos w=2u l=1u
M2918 net880 n2712 VDD VDD pmos w=2u l=1u
M2919 n2812 net881 VDD VDD pmos w=2u l=1u
M2920 net883 net880 VDD VDD pmos w=2u l=1u
M2921 n2711 n2818 VDD VDD pmos w=2u l=1u
M2922 n2711 n2818 VSS VSS nmos w=1u l=1u
M2923 n2811 n2820 net884 VSS nmos w=1u l=1u
M2924 net884 n2819 VSS VSS nmos w=1u l=1u
M2925 n2811 n2820 VDD VDD pmos w=2u l=1u
M2926 n2811 n2819 VDD VDD pmos w=2u l=1u
M2927 net885 n2712 VSS VSS nmos w=1u l=1u
M2928 net886 n2818 VSS VSS nmos w=1u l=1u
M2929 n2820 net887 VSS VSS nmos w=1u l=1u
M2930 net887 n2712 net888 VSS nmos w=1u l=1u
M2931 net887 net885 net886 VSS nmos w=1u l=1u
M2932 net888 net886 VSS VSS nmos w=1u l=1u
M2933 net887 net885 net889 VDD pmos w=2u l=1u
M2934 net885 n2712 VDD VDD pmos w=2u l=1u
M2935 net886 n2712 net887 VDD pmos w=2u l=1u
M2936 net886 n2818 VDD VDD pmos w=2u l=1u
M2937 n2820 net887 VDD VDD pmos w=2u l=1u
M2938 net889 net886 VDD VDD pmos w=2u l=1u
M2939 n2712 N409 net890 VSS nmos w=1u l=1u
M2940 net890 N222 VSS VSS nmos w=1u l=1u
M2941 n2712 N409 VDD VDD pmos w=2u l=1u
M2942 n2712 N222 VDD VDD pmos w=2u l=1u
M2943 n2818 n2709 net891 VSS nmos w=1u l=1u
M2944 net891 n2821 VSS VSS nmos w=1u l=1u
M2945 n2818 n2709 VDD VDD pmos w=2u l=1u
M2946 n2818 n2821 VDD VDD pmos w=2u l=1u
M2947 n2709 n2823 net892 VSS nmos w=1u l=1u
M2948 net892 n2822 VSS VSS nmos w=1u l=1u
M2949 n2709 n2823 VDD VDD pmos w=2u l=1u
M2950 n2709 n2822 VDD VDD pmos w=2u l=1u
M2951 n2823 n2825 net893 VSS nmos w=1u l=1u
M2952 net893 n2824 VSS VSS nmos w=1u l=1u
M2953 n2823 n2825 VDD VDD pmos w=2u l=1u
M2954 n2823 n2824 VDD VDD pmos w=2u l=1u
M2955 n2821 n2824 net894 VSS nmos w=1u l=1u
M2956 net894 n2826 VSS VSS nmos w=1u l=1u
M2957 n2821 n2824 VDD VDD pmos w=2u l=1u
M2958 n2821 n2826 VDD VDD pmos w=2u l=1u
M2959 n2824 n2828 net895 VSS nmos w=1u l=1u
M2960 net895 n2827 VSS VSS nmos w=1u l=1u
M2961 n2824 n2828 VDD VDD pmos w=2u l=1u
M2962 n2824 n2827 VDD VDD pmos w=2u l=1u
M2963 n2826 n2822 VSS VSS nmos w=1u l=1u
M2964 n2826 n2829 VSS VSS nmos w=1u l=1u
M2965 n2826 n2822 net896 VDD pmos w=2u l=1u
M2966 net896 n2829 VDD VDD pmos w=2u l=1u
M2967 n2822 net897 VSS VSS nmos w=1u l=1u
M2968 net898 n2830 VSS VSS nmos w=1u l=1u
M2969 net897 n2724 net898 VSS nmos w=1u l=1u
M2970 net897 n2830 VDD VDD pmos w=2u l=1u
M2971 net897 n2724 VDD VDD pmos w=2u l=1u
M2972 n2822 net897 VDD VDD pmos w=2u l=1u
M2973 n2830 N392 net899 VSS nmos w=1u l=1u
M2974 net899 n2831 VSS VSS nmos w=1u l=1u
M2975 n2830 N392 VDD VDD pmos w=2u l=1u
M2976 n2830 n2831 VDD VDD pmos w=2u l=1u
M2977 n2831 n2833 VSS VSS nmos w=1u l=1u
M2978 n2831 n2832 VSS VSS nmos w=1u l=1u
M2979 n2831 n2833 net900 VDD pmos w=2u l=1u
M2980 net900 n2832 VDD VDD pmos w=2u l=1u
M2981 n2833 n2835 VSS VSS nmos w=1u l=1u
M2982 n2833 n2834 VSS VSS nmos w=1u l=1u
M2983 n2833 n2835 net901 VDD pmos w=2u l=1u
M2984 net901 n2834 VDD VDD pmos w=2u l=1u
M2985 n2835 n2270 net902 VSS nmos w=1u l=1u
M2986 net902 n2836 VSS VSS nmos w=1u l=1u
M2987 n2835 n2270 VDD VDD pmos w=2u l=1u
M2988 n2835 n2836 VDD VDD pmos w=2u l=1u
M2989 n2836 n2837 net903 VSS nmos w=1u l=1u
M2990 net903 N239 VSS VSS nmos w=1u l=1u
M2991 n2836 n2837 VDD VDD pmos w=2u l=1u
M2992 n2836 N239 VDD VDD pmos w=2u l=1u
M2993 n2834 n2727 VDD VDD pmos w=2u l=1u
M2994 n2834 n2727 VSS VSS nmos w=1u l=1u
M2995 n2832 n2727 VSS VSS nmos w=1u l=1u
M2996 n2832 N375 VSS VSS nmos w=1u l=1u
M2997 n2832 n2727 net904 VDD pmos w=2u l=1u
M2998 net904 N375 VDD VDD pmos w=2u l=1u
M2999 n2724 n2839 net905 VSS nmos w=1u l=1u
M3000 net905 n2838 VSS VSS nmos w=1u l=1u
M3001 n2724 n2839 VDD VDD pmos w=2u l=1u
M3002 n2724 n2838 VDD VDD pmos w=2u l=1u
M3003 n2839 N239 net906 VSS nmos w=1u l=1u
M3004 net906 N392 VSS VSS nmos w=1u l=1u
M3005 n2839 N239 VDD VDD pmos w=2u l=1u
M3006 n2839 N392 VDD VDD pmos w=2u l=1u
M3007 net907 n2726 VSS VSS nmos w=1u l=1u
M3008 net908 n2727 VSS VSS nmos w=1u l=1u
M3009 n2838 net909 VSS VSS nmos w=1u l=1u
M3010 net909 n2726 net910 VSS nmos w=1u l=1u
M3011 net909 net907 net908 VSS nmos w=1u l=1u
M3012 net910 net908 VSS VSS nmos w=1u l=1u
M3013 net909 net907 net911 VDD pmos w=2u l=1u
M3014 net907 n2726 VDD VDD pmos w=2u l=1u
M3015 net908 n2726 net909 VDD pmos w=2u l=1u
M3016 net908 n2727 VDD VDD pmos w=2u l=1u
M3017 n2838 net909 VDD VDD pmos w=2u l=1u
M3018 net911 net908 VDD VDD pmos w=2u l=1u
M3019 n2726 N256 net912 VSS nmos w=1u l=1u
M3020 net912 N375 VSS VSS nmos w=1u l=1u
M3021 n2726 N256 VDD VDD pmos w=2u l=1u
M3022 n2726 N375 VDD VDD pmos w=2u l=1u
M3023 n2727 n2841 net913 VSS nmos w=1u l=1u
M3024 net913 n2840 VSS VSS nmos w=1u l=1u
M3025 n2727 n2841 VDD VDD pmos w=2u l=1u
M3026 n2727 n2840 VDD VDD pmos w=2u l=1u
M3027 n2841 n2843 net914 VSS nmos w=1u l=1u
M3028 net914 n2842 VSS VSS nmos w=1u l=1u
M3029 n2841 n2843 VDD VDD pmos w=2u l=1u
M3030 n2841 n2842 VDD VDD pmos w=2u l=1u
M3031 n2829 n2825 VDD VDD pmos w=2u l=1u
M3032 n2829 n2825 VSS VSS nmos w=1u l=1u
M3033 n2819 n2845 VSS VSS nmos w=1u l=1u
M3034 n2819 n2844 VSS VSS nmos w=1u l=1u
M3035 n2819 n2845 net915 VDD pmos w=2u l=1u
M3036 net915 n2844 VDD VDD pmos w=2u l=1u
M3037 n2845 n2816 VSS VSS nmos w=1u l=1u
M3038 n2845 n2817 VSS VSS nmos w=1u l=1u
M3039 n2845 n2816 net916 VDD pmos w=2u l=1u
M3040 net916 n2817 VDD VDD pmos w=2u l=1u
M3041 n2844 n2815 VDD VDD pmos w=2u l=1u
M3042 n2844 n2815 VSS VSS nmos w=1u l=1u
M3043 n2809 n2847 VSS VSS nmos w=1u l=1u
M3044 n2809 n2846 VSS VSS nmos w=1u l=1u
M3045 n2809 n2847 net917 VDD pmos w=2u l=1u
M3046 net917 n2846 VDD VDD pmos w=2u l=1u
M3047 n2847 n2806 VSS VSS nmos w=1u l=1u
M3048 n2847 n2807 VSS VSS nmos w=1u l=1u
M3049 n2847 n2806 net918 VDD pmos w=2u l=1u
M3050 net918 n2807 VDD VDD pmos w=2u l=1u
M3051 n2846 n2805 VDD VDD pmos w=2u l=1u
M3052 n2846 n2805 VSS VSS nmos w=1u l=1u
M3053 n2799 n2849 VSS VSS nmos w=1u l=1u
M3054 n2799 n2848 VSS VSS nmos w=1u l=1u
M3055 n2799 n2849 net919 VDD pmos w=2u l=1u
M3056 net919 n2848 VDD VDD pmos w=2u l=1u
M3057 n2849 n2796 VSS VSS nmos w=1u l=1u
M3058 n2849 n2797 VSS VSS nmos w=1u l=1u
M3059 n2849 n2796 net920 VDD pmos w=2u l=1u
M3060 net920 n2797 VDD VDD pmos w=2u l=1u
M3061 n2848 n2795 VDD VDD pmos w=2u l=1u
M3062 n2848 n2795 VSS VSS nmos w=1u l=1u
M3063 n2789 n2851 VSS VSS nmos w=1u l=1u
M3064 n2789 n2850 VSS VSS nmos w=1u l=1u
M3065 n2789 n2851 net921 VDD pmos w=2u l=1u
M3066 net921 n2850 VDD VDD pmos w=2u l=1u
M3067 n2851 n2786 VSS VSS nmos w=1u l=1u
M3068 n2851 n2787 VSS VSS nmos w=1u l=1u
M3069 n2851 n2786 net922 VDD pmos w=2u l=1u
M3070 net922 n2787 VDD VDD pmos w=2u l=1u
M3071 n2850 n2785 VDD VDD pmos w=2u l=1u
M3072 n2850 n2785 VSS VSS nmos w=1u l=1u
M3073 n2779 n2853 VSS VSS nmos w=1u l=1u
M3074 n2779 n2852 VSS VSS nmos w=1u l=1u
M3075 n2779 n2853 net923 VDD pmos w=2u l=1u
M3076 net923 n2852 VDD VDD pmos w=2u l=1u
M3077 n2853 n2776 VSS VSS nmos w=1u l=1u
M3078 n2853 n2777 VSS VSS nmos w=1u l=1u
M3079 n2853 n2776 net924 VDD pmos w=2u l=1u
M3080 net924 n2777 VDD VDD pmos w=2u l=1u
M3081 n2852 n2775 VDD VDD pmos w=2u l=1u
M3082 n2852 n2775 VSS VSS nmos w=1u l=1u
M3083 n2769 n2855 VSS VSS nmos w=1u l=1u
M3084 n2769 n2854 VSS VSS nmos w=1u l=1u
M3085 n2769 n2855 net925 VDD pmos w=2u l=1u
M3086 net925 n2854 VDD VDD pmos w=2u l=1u
M3087 n2855 n2766 VSS VSS nmos w=1u l=1u
M3088 n2855 n2767 VSS VSS nmos w=1u l=1u
M3089 n2855 n2766 net926 VDD pmos w=2u l=1u
M3090 net926 n2767 VDD VDD pmos w=2u l=1u
M3091 n2854 n2765 VDD VDD pmos w=2u l=1u
M3092 n2854 n2765 VSS VSS nmos w=1u l=1u
M3093 n2759 n2857 VSS VSS nmos w=1u l=1u
M3094 n2759 n2856 VSS VSS nmos w=1u l=1u
M3095 n2759 n2857 net927 VDD pmos w=2u l=1u
M3096 net927 n2856 VDD VDD pmos w=2u l=1u
M3097 n2857 n2756 VSS VSS nmos w=1u l=1u
M3098 n2857 n2757 VSS VSS nmos w=1u l=1u
M3099 n2857 n2756 net928 VDD pmos w=2u l=1u
M3100 net928 n2757 VDD VDD pmos w=2u l=1u
M3101 n2856 n2755 VDD VDD pmos w=2u l=1u
M3102 n2856 n2755 VSS VSS nmos w=1u l=1u
M3103 n2644 N528 net929 VSS nmos w=1u l=1u
M3104 net929 N103 VSS VSS nmos w=1u l=1u
M3105 n2644 N528 VDD VDD pmos w=2u l=1u
M3106 n2644 N103 VDD VDD pmos w=2u l=1u
M3107 N6190 n2858 net930 VSS nmos w=1u l=1u
M3108 net930 n2744 VSS VSS nmos w=1u l=1u
M3109 N6190 n2858 VDD VDD pmos w=2u l=1u
M3110 N6190 n2744 VDD VDD pmos w=2u l=1u
M3111 n2858 net931 VSS VSS nmos w=1u l=1u
M3112 net931 n2859 VSS VSS nmos w=1u l=1u
M3113 net931 n2860 VSS VSS nmos w=1u l=1u
M3114 net931 n2860 net932 VDD pmos w=2u l=1u
M3115 n2858 net931 VDD VDD pmos w=2u l=1u
M3116 net932 n2859 VDD VDD pmos w=2u l=1u
M3117 n2744 n2860 net933 VSS nmos w=1u l=1u
M3118 net933 n2859 VSS VSS nmos w=1u l=1u
M3119 n2744 n2860 VDD VDD pmos w=2u l=1u
M3120 n2744 n2859 VDD VDD pmos w=2u l=1u
M3121 n2860 n2862 net934 VSS nmos w=1u l=1u
M3122 net934 n2861 VSS VSS nmos w=1u l=1u
M3123 n2860 n2862 VDD VDD pmos w=2u l=1u
M3124 n2860 n2861 VDD VDD pmos w=2u l=1u
M3125 n2861 n2864 net935 VSS nmos w=1u l=1u
M3126 net935 n2863 VSS VSS nmos w=1u l=1u
M3127 n2861 n2864 VDD VDD pmos w=2u l=1u
M3128 n2861 n2863 VDD VDD pmos w=2u l=1u
M3129 net936 n2746 VSS VSS nmos w=1u l=1u
M3130 net937 n2745 VSS VSS nmos w=1u l=1u
M3131 n2859 net938 VSS VSS nmos w=1u l=1u
M3132 net938 n2746 net939 VSS nmos w=1u l=1u
M3133 net938 net936 net937 VSS nmos w=1u l=1u
M3134 net939 net937 VSS VSS nmos w=1u l=1u
M3135 net938 net936 net940 VDD pmos w=2u l=1u
M3136 net936 n2746 VDD VDD pmos w=2u l=1u
M3137 net937 n2746 net938 VDD pmos w=2u l=1u
M3138 net937 n2745 VDD VDD pmos w=2u l=1u
M3139 n2859 net938 VDD VDD pmos w=2u l=1u
M3140 net940 net937 VDD VDD pmos w=2u l=1u
M3141 n2746 n2866 net941 VSS nmos w=1u l=1u
M3142 net941 n2865 VSS VSS nmos w=1u l=1u
M3143 n2746 n2866 VDD VDD pmos w=2u l=1u
M3144 n2746 n2865 VDD VDD pmos w=2u l=1u
M3145 n2865 n2868 net942 VSS nmos w=1u l=1u
M3146 net942 n2867 VSS VSS nmos w=1u l=1u
M3147 n2865 n2868 VDD VDD pmos w=2u l=1u
M3148 n2865 n2867 VDD VDD pmos w=2u l=1u
M3149 net943 n2749 VSS VSS nmos w=1u l=1u
M3150 net944 n2750 VSS VSS nmos w=1u l=1u
M3151 n2745 net945 VSS VSS nmos w=1u l=1u
M3152 net945 n2749 net946 VSS nmos w=1u l=1u
M3153 net945 net943 net944 VSS nmos w=1u l=1u
M3154 net946 net944 VSS VSS nmos w=1u l=1u
M3155 net945 net943 net947 VDD pmos w=2u l=1u
M3156 net943 n2749 VDD VDD pmos w=2u l=1u
M3157 net944 n2749 net945 VDD pmos w=2u l=1u
M3158 net944 n2750 VDD VDD pmos w=2u l=1u
M3159 n2745 net945 VDD VDD pmos w=2u l=1u
M3160 net947 net944 VDD VDD pmos w=2u l=1u
M3161 n2749 net948 VSS VSS nmos w=1u l=1u
M3162 net949 n2748 VSS VSS nmos w=1u l=1u
M3163 net948 n2869 net949 VSS nmos w=1u l=1u
M3164 net948 n2748 VDD VDD pmos w=2u l=1u
M3165 net948 n2869 VDD VDD pmos w=2u l=1u
M3166 n2749 net948 VDD VDD pmos w=2u l=1u
M3167 n2748 n2871 net950 VSS nmos w=1u l=1u
M3168 net950 n2870 VSS VSS nmos w=1u l=1u
M3169 n2748 n2871 VDD VDD pmos w=2u l=1u
M3170 n2748 n2870 VDD VDD pmos w=2u l=1u
M3171 n2871 n2873 net951 VSS nmos w=1u l=1u
M3172 net951 n2872 VSS VSS nmos w=1u l=1u
M3173 n2871 n2873 VDD VDD pmos w=2u l=1u
M3174 n2871 n2872 VDD VDD pmos w=2u l=1u
M3175 n2872 net952 VSS VSS nmos w=1u l=1u
M3176 net952 n2874 VSS VSS nmos w=1u l=1u
M3177 net952 n2875 VSS VSS nmos w=1u l=1u
M3178 net952 n2875 net953 VDD pmos w=2u l=1u
M3179 n2872 net952 VDD VDD pmos w=2u l=1u
M3180 net953 n2874 VDD VDD pmos w=2u l=1u
M3181 net954 n2756 VSS VSS nmos w=1u l=1u
M3182 net955 n2757 VSS VSS nmos w=1u l=1u
M3183 n2870 net956 VSS VSS nmos w=1u l=1u
M3184 net956 n2756 net957 VSS nmos w=1u l=1u
M3185 net956 net954 net955 VSS nmos w=1u l=1u
M3186 net957 net955 VSS VSS nmos w=1u l=1u
M3187 net956 net954 net958 VDD pmos w=2u l=1u
M3188 net954 n2756 VDD VDD pmos w=2u l=1u
M3189 net955 n2756 net956 VDD pmos w=2u l=1u
M3190 net955 n2757 VDD VDD pmos w=2u l=1u
M3191 n2870 net956 VDD VDD pmos w=2u l=1u
M3192 net958 net955 VDD VDD pmos w=2u l=1u
M3193 n2757 n2876 VDD VDD pmos w=2u l=1u
M3194 n2757 n2876 VSS VSS nmos w=1u l=1u
M3195 n2869 n2878 net959 VSS nmos w=1u l=1u
M3196 net959 n2877 VSS VSS nmos w=1u l=1u
M3197 n2869 n2878 VDD VDD pmos w=2u l=1u
M3198 n2869 n2877 VDD VDD pmos w=2u l=1u
M3199 net960 n2876 VSS VSS nmos w=1u l=1u
M3200 net961 n2756 VSS VSS nmos w=1u l=1u
M3201 n2878 net962 VSS VSS nmos w=1u l=1u
M3202 net962 n2876 net963 VSS nmos w=1u l=1u
M3203 net962 net960 net961 VSS nmos w=1u l=1u
M3204 net963 net961 VSS VSS nmos w=1u l=1u
M3205 net962 net960 net964 VDD pmos w=2u l=1u
M3206 net960 n2876 VDD VDD pmos w=2u l=1u
M3207 net961 n2876 net962 VDD pmos w=2u l=1u
M3208 net961 n2756 VDD VDD pmos w=2u l=1u
M3209 n2878 net962 VDD VDD pmos w=2u l=1u
M3210 net964 net961 VDD VDD pmos w=2u l=1u
M3211 n2876 N511 net965 VSS nmos w=1u l=1u
M3212 net965 N103 VSS VSS nmos w=1u l=1u
M3213 n2876 N511 VDD VDD pmos w=2u l=1u
M3214 n2876 N103 VDD VDD pmos w=2u l=1u
M3215 n2756 n2755 net966 VSS nmos w=1u l=1u
M3216 net966 n2879 VSS VSS nmos w=1u l=1u
M3217 n2756 n2755 VDD VDD pmos w=2u l=1u
M3218 n2756 n2879 VDD VDD pmos w=2u l=1u
M3219 n2755 n2881 net967 VSS nmos w=1u l=1u
M3220 net967 n2880 VSS VSS nmos w=1u l=1u
M3221 n2755 n2881 VDD VDD pmos w=2u l=1u
M3222 n2755 n2880 VDD VDD pmos w=2u l=1u
M3223 n2881 n2883 net968 VSS nmos w=1u l=1u
M3224 net968 n2882 VSS VSS nmos w=1u l=1u
M3225 n2881 n2883 VDD VDD pmos w=2u l=1u
M3226 n2881 n2882 VDD VDD pmos w=2u l=1u
M3227 n2882 net969 VSS VSS nmos w=1u l=1u
M3228 net969 n2884 VSS VSS nmos w=1u l=1u
M3229 net969 n2885 VSS VSS nmos w=1u l=1u
M3230 net969 n2885 net970 VDD pmos w=2u l=1u
M3231 n2882 net969 VDD VDD pmos w=2u l=1u
M3232 net970 n2884 VDD VDD pmos w=2u l=1u
M3233 net971 n2766 VSS VSS nmos w=1u l=1u
M3234 net972 n2767 VSS VSS nmos w=1u l=1u
M3235 n2880 net973 VSS VSS nmos w=1u l=1u
M3236 net973 n2766 net974 VSS nmos w=1u l=1u
M3237 net973 net971 net972 VSS nmos w=1u l=1u
M3238 net974 net972 VSS VSS nmos w=1u l=1u
M3239 net973 net971 net975 VDD pmos w=2u l=1u
M3240 net971 n2766 VDD VDD pmos w=2u l=1u
M3241 net972 n2766 net973 VDD pmos w=2u l=1u
M3242 net972 n2767 VDD VDD pmos w=2u l=1u
M3243 n2880 net973 VDD VDD pmos w=2u l=1u
M3244 net975 net972 VDD VDD pmos w=2u l=1u
M3245 n2767 n2886 VDD VDD pmos w=2u l=1u
M3246 n2767 n2886 VSS VSS nmos w=1u l=1u
M3247 n2879 n2888 net976 VSS nmos w=1u l=1u
M3248 net976 n2887 VSS VSS nmos w=1u l=1u
M3249 n2879 n2888 VDD VDD pmos w=2u l=1u
M3250 n2879 n2887 VDD VDD pmos w=2u l=1u
M3251 net977 n2886 VSS VSS nmos w=1u l=1u
M3252 net978 n2766 VSS VSS nmos w=1u l=1u
M3253 n2888 net979 VSS VSS nmos w=1u l=1u
M3254 net979 n2886 net980 VSS nmos w=1u l=1u
M3255 net979 net977 net978 VSS nmos w=1u l=1u
M3256 net980 net978 VSS VSS nmos w=1u l=1u
M3257 net979 net977 net981 VDD pmos w=2u l=1u
M3258 net977 n2886 VDD VDD pmos w=2u l=1u
M3259 net978 n2886 net979 VDD pmos w=2u l=1u
M3260 net978 n2766 VDD VDD pmos w=2u l=1u
M3261 n2888 net979 VDD VDD pmos w=2u l=1u
M3262 net981 net978 VDD VDD pmos w=2u l=1u
M3263 n2886 N494 net982 VSS nmos w=1u l=1u
M3264 net982 N120 VSS VSS nmos w=1u l=1u
M3265 n2886 N494 VDD VDD pmos w=2u l=1u
M3266 n2886 N120 VDD VDD pmos w=2u l=1u
M3267 n2766 n2765 net983 VSS nmos w=1u l=1u
M3268 net983 n2889 VSS VSS nmos w=1u l=1u
M3269 n2766 n2765 VDD VDD pmos w=2u l=1u
M3270 n2766 n2889 VDD VDD pmos w=2u l=1u
M3271 n2765 n2891 net984 VSS nmos w=1u l=1u
M3272 net984 n2890 VSS VSS nmos w=1u l=1u
M3273 n2765 n2891 VDD VDD pmos w=2u l=1u
M3274 n2765 n2890 VDD VDD pmos w=2u l=1u
M3275 n2891 n2893 net985 VSS nmos w=1u l=1u
M3276 net985 n2892 VSS VSS nmos w=1u l=1u
M3277 n2891 n2893 VDD VDD pmos w=2u l=1u
M3278 n2891 n2892 VDD VDD pmos w=2u l=1u
M3279 n2892 net986 VSS VSS nmos w=1u l=1u
M3280 net986 n2894 VSS VSS nmos w=1u l=1u
M3281 net986 n2895 VSS VSS nmos w=1u l=1u
M3282 net986 n2895 net987 VDD pmos w=2u l=1u
M3283 n2892 net986 VDD VDD pmos w=2u l=1u
M3284 net987 n2894 VDD VDD pmos w=2u l=1u
M3285 net988 n2776 VSS VSS nmos w=1u l=1u
M3286 net989 n2777 VSS VSS nmos w=1u l=1u
M3287 n2890 net990 VSS VSS nmos w=1u l=1u
M3288 net990 n2776 net991 VSS nmos w=1u l=1u
M3289 net990 net988 net989 VSS nmos w=1u l=1u
M3290 net991 net989 VSS VSS nmos w=1u l=1u
M3291 net990 net988 net992 VDD pmos w=2u l=1u
M3292 net988 n2776 VDD VDD pmos w=2u l=1u
M3293 net989 n2776 net990 VDD pmos w=2u l=1u
M3294 net989 n2777 VDD VDD pmos w=2u l=1u
M3295 n2890 net990 VDD VDD pmos w=2u l=1u
M3296 net992 net989 VDD VDD pmos w=2u l=1u
M3297 n2777 n2896 VDD VDD pmos w=2u l=1u
M3298 n2777 n2896 VSS VSS nmos w=1u l=1u
M3299 n2889 n2898 net993 VSS nmos w=1u l=1u
M3300 net993 n2897 VSS VSS nmos w=1u l=1u
M3301 n2889 n2898 VDD VDD pmos w=2u l=1u
M3302 n2889 n2897 VDD VDD pmos w=2u l=1u
M3303 net994 n2896 VSS VSS nmos w=1u l=1u
M3304 net995 n2776 VSS VSS nmos w=1u l=1u
M3305 n2898 net996 VSS VSS nmos w=1u l=1u
M3306 net996 n2896 net997 VSS nmos w=1u l=1u
M3307 net996 net994 net995 VSS nmos w=1u l=1u
M3308 net997 net995 VSS VSS nmos w=1u l=1u
M3309 net996 net994 net998 VDD pmos w=2u l=1u
M3310 net994 n2896 VDD VDD pmos w=2u l=1u
M3311 net995 n2896 net996 VDD pmos w=2u l=1u
M3312 net995 n2776 VDD VDD pmos w=2u l=1u
M3313 n2898 net996 VDD VDD pmos w=2u l=1u
M3314 net998 net995 VDD VDD pmos w=2u l=1u
M3315 n2896 N477 net999 VSS nmos w=1u l=1u
M3316 net999 N137 VSS VSS nmos w=1u l=1u
M3317 n2896 N477 VDD VDD pmos w=2u l=1u
M3318 n2896 N137 VDD VDD pmos w=2u l=1u
M3319 n2776 n2775 net1000 VSS nmos w=1u l=1u
M3320 net1000 n2899 VSS VSS nmos w=1u l=1u
M3321 n2776 n2775 VDD VDD pmos w=2u l=1u
M3322 n2776 n2899 VDD VDD pmos w=2u l=1u
M3323 n2775 n2901 net1001 VSS nmos w=1u l=1u
M3324 net1001 n2900 VSS VSS nmos w=1u l=1u
M3325 n2775 n2901 VDD VDD pmos w=2u l=1u
M3326 n2775 n2900 VDD VDD pmos w=2u l=1u
M3327 n2901 n2903 net1002 VSS nmos w=1u l=1u
M3328 net1002 n2902 VSS VSS nmos w=1u l=1u
M3329 n2901 n2903 VDD VDD pmos w=2u l=1u
M3330 n2901 n2902 VDD VDD pmos w=2u l=1u
M3331 n2902 net1003 VSS VSS nmos w=1u l=1u
M3332 net1003 n2904 VSS VSS nmos w=1u l=1u
M3333 net1003 n2905 VSS VSS nmos w=1u l=1u
M3334 net1003 n2905 net1004 VDD pmos w=2u l=1u
M3335 n2902 net1003 VDD VDD pmos w=2u l=1u
M3336 net1004 n2904 VDD VDD pmos w=2u l=1u
M3337 net1005 n2786 VSS VSS nmos w=1u l=1u
M3338 net1006 n2787 VSS VSS nmos w=1u l=1u
M3339 n2900 net1007 VSS VSS nmos w=1u l=1u
M3340 net1007 n2786 net1008 VSS nmos w=1u l=1u
M3341 net1007 net1005 net1006 VSS nmos w=1u l=1u
M3342 net1008 net1006 VSS VSS nmos w=1u l=1u
M3343 net1007 net1005 net1009 VDD pmos w=2u l=1u
M3344 net1005 n2786 VDD VDD pmos w=2u l=1u
M3345 net1006 n2786 net1007 VDD pmos w=2u l=1u
M3346 net1006 n2787 VDD VDD pmos w=2u l=1u
M3347 n2900 net1007 VDD VDD pmos w=2u l=1u
M3348 net1009 net1006 VDD VDD pmos w=2u l=1u
M3349 n2787 n2906 VDD VDD pmos w=2u l=1u
M3350 n2787 n2906 VSS VSS nmos w=1u l=1u
M3351 n2899 n2908 net1010 VSS nmos w=1u l=1u
M3352 net1010 n2907 VSS VSS nmos w=1u l=1u
M3353 n2899 n2908 VDD VDD pmos w=2u l=1u
M3354 n2899 n2907 VDD VDD pmos w=2u l=1u
M3355 net1011 n2906 VSS VSS nmos w=1u l=1u
M3356 net1012 n2786 VSS VSS nmos w=1u l=1u
M3357 n2908 net1013 VSS VSS nmos w=1u l=1u
M3358 net1013 n2906 net1014 VSS nmos w=1u l=1u
M3359 net1013 net1011 net1012 VSS nmos w=1u l=1u
M3360 net1014 net1012 VSS VSS nmos w=1u l=1u
M3361 net1013 net1011 net1015 VDD pmos w=2u l=1u
M3362 net1011 n2906 VDD VDD pmos w=2u l=1u
M3363 net1012 n2906 net1013 VDD pmos w=2u l=1u
M3364 net1012 n2786 VDD VDD pmos w=2u l=1u
M3365 n2908 net1013 VDD VDD pmos w=2u l=1u
M3366 net1015 net1012 VDD VDD pmos w=2u l=1u
M3367 n2906 N460 net1016 VSS nmos w=1u l=1u
M3368 net1016 N154 VSS VSS nmos w=1u l=1u
M3369 n2906 N460 VDD VDD pmos w=2u l=1u
M3370 n2906 N154 VDD VDD pmos w=2u l=1u
M3371 n2786 n2785 net1017 VSS nmos w=1u l=1u
M3372 net1017 n2909 VSS VSS nmos w=1u l=1u
M3373 n2786 n2785 VDD VDD pmos w=2u l=1u
M3374 n2786 n2909 VDD VDD pmos w=2u l=1u
M3375 n2785 n2911 net1018 VSS nmos w=1u l=1u
M3376 net1018 n2910 VSS VSS nmos w=1u l=1u
M3377 n2785 n2911 VDD VDD pmos w=2u l=1u
M3378 n2785 n2910 VDD VDD pmos w=2u l=1u
M3379 n2911 n2913 net1019 VSS nmos w=1u l=1u
M3380 net1019 n2912 VSS VSS nmos w=1u l=1u
M3381 n2911 n2913 VDD VDD pmos w=2u l=1u
M3382 n2911 n2912 VDD VDD pmos w=2u l=1u
M3383 n2912 net1020 VSS VSS nmos w=1u l=1u
M3384 net1020 n2914 VSS VSS nmos w=1u l=1u
M3385 net1020 n2915 VSS VSS nmos w=1u l=1u
M3386 net1020 n2915 net1021 VDD pmos w=2u l=1u
M3387 n2912 net1020 VDD VDD pmos w=2u l=1u
M3388 net1021 n2914 VDD VDD pmos w=2u l=1u
M3389 net1022 n2796 VSS VSS nmos w=1u l=1u
M3390 net1023 n2797 VSS VSS nmos w=1u l=1u
M3391 n2910 net1024 VSS VSS nmos w=1u l=1u
M3392 net1024 n2796 net1025 VSS nmos w=1u l=1u
M3393 net1024 net1022 net1023 VSS nmos w=1u l=1u
M3394 net1025 net1023 VSS VSS nmos w=1u l=1u
M3395 net1024 net1022 net1026 VDD pmos w=2u l=1u
M3396 net1022 n2796 VDD VDD pmos w=2u l=1u
M3397 net1023 n2796 net1024 VDD pmos w=2u l=1u
M3398 net1023 n2797 VDD VDD pmos w=2u l=1u
M3399 n2910 net1024 VDD VDD pmos w=2u l=1u
M3400 net1026 net1023 VDD VDD pmos w=2u l=1u
M3401 n2797 n2916 VDD VDD pmos w=2u l=1u
M3402 n2797 n2916 VSS VSS nmos w=1u l=1u
M3403 n2909 n2918 net1027 VSS nmos w=1u l=1u
M3404 net1027 n2917 VSS VSS nmos w=1u l=1u
M3405 n2909 n2918 VDD VDD pmos w=2u l=1u
M3406 n2909 n2917 VDD VDD pmos w=2u l=1u
M3407 net1028 n2916 VSS VSS nmos w=1u l=1u
M3408 net1029 n2796 VSS VSS nmos w=1u l=1u
M3409 n2918 net1030 VSS VSS nmos w=1u l=1u
M3410 net1030 n2916 net1031 VSS nmos w=1u l=1u
M3411 net1030 net1028 net1029 VSS nmos w=1u l=1u
M3412 net1031 net1029 VSS VSS nmos w=1u l=1u
M3413 net1030 net1028 net1032 VDD pmos w=2u l=1u
M3414 net1028 n2916 VDD VDD pmos w=2u l=1u
M3415 net1029 n2916 net1030 VDD pmos w=2u l=1u
M3416 net1029 n2796 VDD VDD pmos w=2u l=1u
M3417 n2918 net1030 VDD VDD pmos w=2u l=1u
M3418 net1032 net1029 VDD VDD pmos w=2u l=1u
M3419 n2916 N443 net1033 VSS nmos w=1u l=1u
M3420 net1033 N171 VSS VSS nmos w=1u l=1u
M3421 n2916 N443 VDD VDD pmos w=2u l=1u
M3422 n2916 N171 VDD VDD pmos w=2u l=1u
M3423 n2796 n2795 net1034 VSS nmos w=1u l=1u
M3424 net1034 n2919 VSS VSS nmos w=1u l=1u
M3425 n2796 n2795 VDD VDD pmos w=2u l=1u
M3426 n2796 n2919 VDD VDD pmos w=2u l=1u
M3427 n2795 n2921 net1035 VSS nmos w=1u l=1u
M3428 net1035 n2920 VSS VSS nmos w=1u l=1u
M3429 n2795 n2921 VDD VDD pmos w=2u l=1u
M3430 n2795 n2920 VDD VDD pmos w=2u l=1u
M3431 n2921 n2923 net1036 VSS nmos w=1u l=1u
M3432 net1036 n2922 VSS VSS nmos w=1u l=1u
M3433 n2921 n2923 VDD VDD pmos w=2u l=1u
M3434 n2921 n2922 VDD VDD pmos w=2u l=1u
M3435 n2922 net1037 VSS VSS nmos w=1u l=1u
M3436 net1037 n2924 VSS VSS nmos w=1u l=1u
M3437 net1037 n2925 VSS VSS nmos w=1u l=1u
M3438 net1037 n2925 net1038 VDD pmos w=2u l=1u
M3439 n2922 net1037 VDD VDD pmos w=2u l=1u
M3440 net1038 n2924 VDD VDD pmos w=2u l=1u
M3441 net1039 n2806 VSS VSS nmos w=1u l=1u
M3442 net1040 n2807 VSS VSS nmos w=1u l=1u
M3443 n2920 net1041 VSS VSS nmos w=1u l=1u
M3444 net1041 n2806 net1042 VSS nmos w=1u l=1u
M3445 net1041 net1039 net1040 VSS nmos w=1u l=1u
M3446 net1042 net1040 VSS VSS nmos w=1u l=1u
M3447 net1041 net1039 net1043 VDD pmos w=2u l=1u
M3448 net1039 n2806 VDD VDD pmos w=2u l=1u
M3449 net1040 n2806 net1041 VDD pmos w=2u l=1u
M3450 net1040 n2807 VDD VDD pmos w=2u l=1u
M3451 n2920 net1041 VDD VDD pmos w=2u l=1u
M3452 net1043 net1040 VDD VDD pmos w=2u l=1u
M3453 n2807 n2926 VDD VDD pmos w=2u l=1u
M3454 n2807 n2926 VSS VSS nmos w=1u l=1u
M3455 n2919 n2928 net1044 VSS nmos w=1u l=1u
M3456 net1044 n2927 VSS VSS nmos w=1u l=1u
M3457 n2919 n2928 VDD VDD pmos w=2u l=1u
M3458 n2919 n2927 VDD VDD pmos w=2u l=1u
M3459 net1045 n2926 VSS VSS nmos w=1u l=1u
M3460 net1046 n2806 VSS VSS nmos w=1u l=1u
M3461 n2928 net1047 VSS VSS nmos w=1u l=1u
M3462 net1047 n2926 net1048 VSS nmos w=1u l=1u
M3463 net1047 net1045 net1046 VSS nmos w=1u l=1u
M3464 net1048 net1046 VSS VSS nmos w=1u l=1u
M3465 net1047 net1045 net1049 VDD pmos w=2u l=1u
M3466 net1045 n2926 VDD VDD pmos w=2u l=1u
M3467 net1046 n2926 net1047 VDD pmos w=2u l=1u
M3468 net1046 n2806 VDD VDD pmos w=2u l=1u
M3469 n2928 net1047 VDD VDD pmos w=2u l=1u
M3470 net1049 net1046 VDD VDD pmos w=2u l=1u
M3471 n2926 N426 net1050 VSS nmos w=1u l=1u
M3472 net1050 N188 VSS VSS nmos w=1u l=1u
M3473 n2926 N426 VDD VDD pmos w=2u l=1u
M3474 n2926 N188 VDD VDD pmos w=2u l=1u
M3475 n2806 n2805 net1051 VSS nmos w=1u l=1u
M3476 net1051 n2929 VSS VSS nmos w=1u l=1u
M3477 n2806 n2805 VDD VDD pmos w=2u l=1u
M3478 n2806 n2929 VDD VDD pmos w=2u l=1u
M3479 n2805 n2931 net1052 VSS nmos w=1u l=1u
M3480 net1052 n2930 VSS VSS nmos w=1u l=1u
M3481 n2805 n2931 VDD VDD pmos w=2u l=1u
M3482 n2805 n2930 VDD VDD pmos w=2u l=1u
M3483 n2931 n2933 net1053 VSS nmos w=1u l=1u
M3484 net1053 n2932 VSS VSS nmos w=1u l=1u
M3485 n2931 n2933 VDD VDD pmos w=2u l=1u
M3486 n2931 n2932 VDD VDD pmos w=2u l=1u
M3487 n2932 net1054 VSS VSS nmos w=1u l=1u
M3488 net1054 n2934 VSS VSS nmos w=1u l=1u
M3489 net1054 n2935 VSS VSS nmos w=1u l=1u
M3490 net1054 n2935 net1055 VDD pmos w=2u l=1u
M3491 n2932 net1054 VDD VDD pmos w=2u l=1u
M3492 net1055 n2934 VDD VDD pmos w=2u l=1u
M3493 net1056 n2816 VSS VSS nmos w=1u l=1u
M3494 net1057 n2817 VSS VSS nmos w=1u l=1u
M3495 n2930 net1058 VSS VSS nmos w=1u l=1u
M3496 net1058 n2816 net1059 VSS nmos w=1u l=1u
M3497 net1058 net1056 net1057 VSS nmos w=1u l=1u
M3498 net1059 net1057 VSS VSS nmos w=1u l=1u
M3499 net1058 net1056 net1060 VDD pmos w=2u l=1u
M3500 net1056 n2816 VDD VDD pmos w=2u l=1u
M3501 net1057 n2816 net1058 VDD pmos w=2u l=1u
M3502 net1057 n2817 VDD VDD pmos w=2u l=1u
M3503 n2930 net1058 VDD VDD pmos w=2u l=1u
M3504 net1060 net1057 VDD VDD pmos w=2u l=1u
M3505 n2817 n2936 VDD VDD pmos w=2u l=1u
M3506 n2817 n2936 VSS VSS nmos w=1u l=1u
M3507 n2929 n2938 net1061 VSS nmos w=1u l=1u
M3508 net1061 n2937 VSS VSS nmos w=1u l=1u
M3509 n2929 n2938 VDD VDD pmos w=2u l=1u
M3510 n2929 n2937 VDD VDD pmos w=2u l=1u
M3511 net1062 n2936 VSS VSS nmos w=1u l=1u
M3512 net1063 n2816 VSS VSS nmos w=1u l=1u
M3513 n2938 net1064 VSS VSS nmos w=1u l=1u
M3514 net1064 n2936 net1065 VSS nmos w=1u l=1u
M3515 net1064 net1062 net1063 VSS nmos w=1u l=1u
M3516 net1065 net1063 VSS VSS nmos w=1u l=1u
M3517 net1064 net1062 net1066 VDD pmos w=2u l=1u
M3518 net1062 n2936 VDD VDD pmos w=2u l=1u
M3519 net1063 n2936 net1064 VDD pmos w=2u l=1u
M3520 net1063 n2816 VDD VDD pmos w=2u l=1u
M3521 n2938 net1064 VDD VDD pmos w=2u l=1u
M3522 net1066 net1063 VDD VDD pmos w=2u l=1u
M3523 n2936 N409 net1067 VSS nmos w=1u l=1u
M3524 net1067 N205 VSS VSS nmos w=1u l=1u
M3525 n2936 N409 VDD VDD pmos w=2u l=1u
M3526 n2936 N205 VDD VDD pmos w=2u l=1u
M3527 n2816 n2815 net1068 VSS nmos w=1u l=1u
M3528 net1068 n2939 VSS VSS nmos w=1u l=1u
M3529 n2816 n2815 VDD VDD pmos w=2u l=1u
M3530 n2816 n2939 VDD VDD pmos w=2u l=1u
M3531 n2815 n2941 net1069 VSS nmos w=1u l=1u
M3532 net1069 n2940 VSS VSS nmos w=1u l=1u
M3533 n2815 n2941 VDD VDD pmos w=2u l=1u
M3534 n2815 n2940 VDD VDD pmos w=2u l=1u
M3535 n2941 n2943 net1070 VSS nmos w=1u l=1u
M3536 net1070 n2942 VSS VSS nmos w=1u l=1u
M3537 n2941 n2943 VDD VDD pmos w=2u l=1u
M3538 n2941 n2942 VDD VDD pmos w=2u l=1u
M3539 n2942 n2945 net1071 VSS nmos w=1u l=1u
M3540 net1071 n2944 VSS VSS nmos w=1u l=1u
M3541 n2942 n2945 VDD VDD pmos w=2u l=1u
M3542 n2942 n2944 VDD VDD pmos w=2u l=1u
M3543 net1072 n2827 VSS VSS nmos w=1u l=1u
M3544 net1073 n2828 VSS VSS nmos w=1u l=1u
M3545 n2940 net1074 VSS VSS nmos w=1u l=1u
M3546 net1074 n2827 net1075 VSS nmos w=1u l=1u
M3547 net1074 net1072 net1073 VSS nmos w=1u l=1u
M3548 net1075 net1073 VSS VSS nmos w=1u l=1u
M3549 net1074 net1072 net1076 VDD pmos w=2u l=1u
M3550 net1072 n2827 VDD VDD pmos w=2u l=1u
M3551 net1073 n2827 net1074 VDD pmos w=2u l=1u
M3552 net1073 n2828 VDD VDD pmos w=2u l=1u
M3553 n2940 net1074 VDD VDD pmos w=2u l=1u
M3554 net1076 net1073 VDD VDD pmos w=2u l=1u
M3555 n2827 n2946 VDD VDD pmos w=2u l=1u
M3556 n2827 n2946 VSS VSS nmos w=1u l=1u
M3557 n2939 n2948 net1077 VSS nmos w=1u l=1u
M3558 net1077 n2947 VSS VSS nmos w=1u l=1u
M3559 n2939 n2948 VDD VDD pmos w=2u l=1u
M3560 n2939 n2947 VDD VDD pmos w=2u l=1u
M3561 net1078 n2828 VSS VSS nmos w=1u l=1u
M3562 net1079 n2946 VSS VSS nmos w=1u l=1u
M3563 n2948 net1080 VSS VSS nmos w=1u l=1u
M3564 net1080 n2828 net1081 VSS nmos w=1u l=1u
M3565 net1080 net1078 net1079 VSS nmos w=1u l=1u
M3566 net1081 net1079 VSS VSS nmos w=1u l=1u
M3567 net1080 net1078 net1082 VDD pmos w=2u l=1u
M3568 net1078 n2828 VDD VDD pmos w=2u l=1u
M3569 net1079 n2828 net1080 VDD pmos w=2u l=1u
M3570 net1079 n2946 VDD VDD pmos w=2u l=1u
M3571 n2948 net1080 VDD VDD pmos w=2u l=1u
M3572 net1082 net1079 VDD VDD pmos w=2u l=1u
M3573 n2828 N392 net1083 VSS nmos w=1u l=1u
M3574 net1083 N222 VSS VSS nmos w=1u l=1u
M3575 n2828 N392 VDD VDD pmos w=2u l=1u
M3576 n2828 N222 VDD VDD pmos w=2u l=1u
M3577 n2946 n2825 net1084 VSS nmos w=1u l=1u
M3578 net1084 n2949 VSS VSS nmos w=1u l=1u
M3579 n2946 n2825 VDD VDD pmos w=2u l=1u
M3580 n2946 n2949 VDD VDD pmos w=2u l=1u
M3581 n2825 n2951 net1085 VSS nmos w=1u l=1u
M3582 net1085 n2950 VSS VSS nmos w=1u l=1u
M3583 n2825 n2951 VDD VDD pmos w=2u l=1u
M3584 n2825 n2950 VDD VDD pmos w=2u l=1u
M3585 n2951 n2953 net1086 VSS nmos w=1u l=1u
M3586 net1086 n2952 VSS VSS nmos w=1u l=1u
M3587 n2951 n2953 VDD VDD pmos w=2u l=1u
M3588 n2951 n2952 VDD VDD pmos w=2u l=1u
M3589 n2949 n2952 net1087 VSS nmos w=1u l=1u
M3590 net1087 n2954 VSS VSS nmos w=1u l=1u
M3591 n2949 n2952 VDD VDD pmos w=2u l=1u
M3592 n2949 n2954 VDD VDD pmos w=2u l=1u
M3593 n2952 n2956 net1088 VSS nmos w=1u l=1u
M3594 net1088 n2955 VSS VSS nmos w=1u l=1u
M3595 n2952 n2956 VDD VDD pmos w=2u l=1u
M3596 n2952 n2955 VDD VDD pmos w=2u l=1u
M3597 n2954 n2950 VSS VSS nmos w=1u l=1u
M3598 n2954 n2957 VSS VSS nmos w=1u l=1u
M3599 n2954 n2950 net1089 VDD pmos w=2u l=1u
M3600 net1089 n2957 VDD VDD pmos w=2u l=1u
M3601 n2950 net1090 VSS VSS nmos w=1u l=1u
M3602 net1091 n2958 VSS VSS nmos w=1u l=1u
M3603 net1090 n2840 net1091 VSS nmos w=1u l=1u
M3604 net1090 n2958 VDD VDD pmos w=2u l=1u
M3605 net1090 n2840 VDD VDD pmos w=2u l=1u
M3606 n2950 net1090 VDD VDD pmos w=2u l=1u
M3607 n2958 N375 net1092 VSS nmos w=1u l=1u
M3608 net1092 n2959 VSS VSS nmos w=1u l=1u
M3609 n2958 N375 VDD VDD pmos w=2u l=1u
M3610 n2958 n2959 VDD VDD pmos w=2u l=1u
M3611 n2959 n2961 VSS VSS nmos w=1u l=1u
M3612 n2959 n2960 VSS VSS nmos w=1u l=1u
M3613 n2959 n2961 net1093 VDD pmos w=2u l=1u
M3614 net1093 n2960 VDD VDD pmos w=2u l=1u
M3615 n2961 n2963 VSS VSS nmos w=1u l=1u
M3616 n2961 n2962 VSS VSS nmos w=1u l=1u
M3617 n2961 n2963 net1094 VDD pmos w=2u l=1u
M3618 net1094 n2962 VDD VDD pmos w=2u l=1u
M3619 n2963 n2270 net1095 VSS nmos w=1u l=1u
M3620 net1095 n2964 VSS VSS nmos w=1u l=1u
M3621 n2963 n2270 VDD VDD pmos w=2u l=1u
M3622 n2963 n2964 VDD VDD pmos w=2u l=1u
M3623 n2964 n2965 net1096 VSS nmos w=1u l=1u
M3624 net1096 N239 VSS VSS nmos w=1u l=1u
M3625 n2964 n2965 VDD VDD pmos w=2u l=1u
M3626 n2964 N239 VDD VDD pmos w=2u l=1u
M3627 n2962 n2843 VDD VDD pmos w=2u l=1u
M3628 n2962 n2843 VSS VSS nmos w=1u l=1u
M3629 n2960 n2843 VSS VSS nmos w=1u l=1u
M3630 n2960 N358 VSS VSS nmos w=1u l=1u
M3631 n2960 n2843 net1097 VDD pmos w=2u l=1u
M3632 net1097 N358 VDD VDD pmos w=2u l=1u
M3633 n2840 n2967 net1098 VSS nmos w=1u l=1u
M3634 net1098 n2966 VSS VSS nmos w=1u l=1u
M3635 n2840 n2967 VDD VDD pmos w=2u l=1u
M3636 n2840 n2966 VDD VDD pmos w=2u l=1u
M3637 n2967 N239 net1099 VSS nmos w=1u l=1u
M3638 net1099 N375 VSS VSS nmos w=1u l=1u
M3639 n2967 N239 VDD VDD pmos w=2u l=1u
M3640 n2967 N375 VDD VDD pmos w=2u l=1u
M3641 net1100 n2842 VSS VSS nmos w=1u l=1u
M3642 net1101 n2843 VSS VSS nmos w=1u l=1u
M3643 n2966 net1102 VSS VSS nmos w=1u l=1u
M3644 net1102 n2842 net1103 VSS nmos w=1u l=1u
M3645 net1102 net1100 net1101 VSS nmos w=1u l=1u
M3646 net1103 net1101 VSS VSS nmos w=1u l=1u
M3647 net1102 net1100 net1104 VDD pmos w=2u l=1u
M3648 net1100 n2842 VDD VDD pmos w=2u l=1u
M3649 net1101 n2842 net1102 VDD pmos w=2u l=1u
M3650 net1101 n2843 VDD VDD pmos w=2u l=1u
M3651 n2966 net1102 VDD VDD pmos w=2u l=1u
M3652 net1104 net1101 VDD VDD pmos w=2u l=1u
M3653 n2842 N256 net1105 VSS nmos w=1u l=1u
M3654 net1105 N358 VSS VSS nmos w=1u l=1u
M3655 n2842 N256 VDD VDD pmos w=2u l=1u
M3656 n2842 N358 VDD VDD pmos w=2u l=1u
M3657 n2843 n2969 net1106 VSS nmos w=1u l=1u
M3658 net1106 n2968 VSS VSS nmos w=1u l=1u
M3659 n2843 n2969 VDD VDD pmos w=2u l=1u
M3660 n2843 n2968 VDD VDD pmos w=2u l=1u
M3661 n2969 n2971 net1107 VSS nmos w=1u l=1u
M3662 net1107 n2970 VSS VSS nmos w=1u l=1u
M3663 n2969 n2971 VDD VDD pmos w=2u l=1u
M3664 n2969 n2970 VDD VDD pmos w=2u l=1u
M3665 n2957 n2953 VDD VDD pmos w=2u l=1u
M3666 n2957 n2953 VSS VSS nmos w=1u l=1u
M3667 n2947 n2973 VSS VSS nmos w=1u l=1u
M3668 n2947 n2972 VSS VSS nmos w=1u l=1u
M3669 n2947 n2973 net1108 VDD pmos w=2u l=1u
M3670 net1108 n2972 VDD VDD pmos w=2u l=1u
M3671 n2973 net1109 VSS VSS nmos w=1u l=1u
M3672 net1110 n2944 VSS VSS nmos w=1u l=1u
M3673 net1109 n2945 net1110 VSS nmos w=1u l=1u
M3674 net1109 n2944 VDD VDD pmos w=2u l=1u
M3675 net1109 n2945 VDD VDD pmos w=2u l=1u
M3676 n2973 net1109 VDD VDD pmos w=2u l=1u
M3677 n2972 n2943 VDD VDD pmos w=2u l=1u
M3678 n2972 n2943 VSS VSS nmos w=1u l=1u
M3679 n2937 n2975 VSS VSS nmos w=1u l=1u
M3680 n2937 n2974 VSS VSS nmos w=1u l=1u
M3681 n2937 n2975 net1111 VDD pmos w=2u l=1u
M3682 net1111 n2974 VDD VDD pmos w=2u l=1u
M3683 n2975 n2934 VSS VSS nmos w=1u l=1u
M3684 n2975 n2935 VSS VSS nmos w=1u l=1u
M3685 n2975 n2934 net1112 VDD pmos w=2u l=1u
M3686 net1112 n2935 VDD VDD pmos w=2u l=1u
M3687 n2974 n2933 VDD VDD pmos w=2u l=1u
M3688 n2974 n2933 VSS VSS nmos w=1u l=1u
M3689 n2927 n2977 VSS VSS nmos w=1u l=1u
M3690 n2927 n2976 VSS VSS nmos w=1u l=1u
M3691 n2927 n2977 net1113 VDD pmos w=2u l=1u
M3692 net1113 n2976 VDD VDD pmos w=2u l=1u
M3693 n2977 n2924 VSS VSS nmos w=1u l=1u
M3694 n2977 n2925 VSS VSS nmos w=1u l=1u
M3695 n2977 n2924 net1114 VDD pmos w=2u l=1u
M3696 net1114 n2925 VDD VDD pmos w=2u l=1u
M3697 n2976 n2923 VDD VDD pmos w=2u l=1u
M3698 n2976 n2923 VSS VSS nmos w=1u l=1u
M3699 n2917 n2979 VSS VSS nmos w=1u l=1u
M3700 n2917 n2978 VSS VSS nmos w=1u l=1u
M3701 n2917 n2979 net1115 VDD pmos w=2u l=1u
M3702 net1115 n2978 VDD VDD pmos w=2u l=1u
M3703 n2979 n2914 VSS VSS nmos w=1u l=1u
M3704 n2979 n2915 VSS VSS nmos w=1u l=1u
M3705 n2979 n2914 net1116 VDD pmos w=2u l=1u
M3706 net1116 n2915 VDD VDD pmos w=2u l=1u
M3707 n2978 n2913 VDD VDD pmos w=2u l=1u
M3708 n2978 n2913 VSS VSS nmos w=1u l=1u
M3709 n2907 n2981 VSS VSS nmos w=1u l=1u
M3710 n2907 n2980 VSS VSS nmos w=1u l=1u
M3711 n2907 n2981 net1117 VDD pmos w=2u l=1u
M3712 net1117 n2980 VDD VDD pmos w=2u l=1u
M3713 n2981 n2904 VSS VSS nmos w=1u l=1u
M3714 n2981 n2905 VSS VSS nmos w=1u l=1u
M3715 n2981 n2904 net1118 VDD pmos w=2u l=1u
M3716 net1118 n2905 VDD VDD pmos w=2u l=1u
M3717 n2980 n2903 VDD VDD pmos w=2u l=1u
M3718 n2980 n2903 VSS VSS nmos w=1u l=1u
M3719 n2897 n2983 VSS VSS nmos w=1u l=1u
M3720 n2897 n2982 VSS VSS nmos w=1u l=1u
M3721 n2897 n2983 net1119 VDD pmos w=2u l=1u
M3722 net1119 n2982 VDD VDD pmos w=2u l=1u
M3723 n2983 n2894 VSS VSS nmos w=1u l=1u
M3724 n2983 n2895 VSS VSS nmos w=1u l=1u
M3725 n2983 n2894 net1120 VDD pmos w=2u l=1u
M3726 net1120 n2895 VDD VDD pmos w=2u l=1u
M3727 n2982 n2893 VDD VDD pmos w=2u l=1u
M3728 n2982 n2893 VSS VSS nmos w=1u l=1u
M3729 n2887 n2985 VSS VSS nmos w=1u l=1u
M3730 n2887 n2984 VSS VSS nmos w=1u l=1u
M3731 n2887 n2985 net1121 VDD pmos w=2u l=1u
M3732 net1121 n2984 VDD VDD pmos w=2u l=1u
M3733 n2985 n2884 VSS VSS nmos w=1u l=1u
M3734 n2985 n2885 VSS VSS nmos w=1u l=1u
M3735 n2985 n2884 net1122 VDD pmos w=2u l=1u
M3736 net1122 n2885 VDD VDD pmos w=2u l=1u
M3737 n2984 n2883 VDD VDD pmos w=2u l=1u
M3738 n2984 n2883 VSS VSS nmos w=1u l=1u
M3739 n2877 n2987 VSS VSS nmos w=1u l=1u
M3740 n2877 n2986 VSS VSS nmos w=1u l=1u
M3741 n2877 n2987 net1123 VDD pmos w=2u l=1u
M3742 net1123 n2986 VDD VDD pmos w=2u l=1u
M3743 n2987 n2874 VSS VSS nmos w=1u l=1u
M3744 n2987 n2875 VSS VSS nmos w=1u l=1u
M3745 n2987 n2874 net1124 VDD pmos w=2u l=1u
M3746 net1124 n2875 VDD VDD pmos w=2u l=1u
M3747 n2986 n2873 VDD VDD pmos w=2u l=1u
M3748 n2986 n2873 VSS VSS nmos w=1u l=1u
M3749 n2750 N528 net1125 VSS nmos w=1u l=1u
M3750 net1125 N86 VSS VSS nmos w=1u l=1u
M3751 n2750 N528 VDD VDD pmos w=2u l=1u
M3752 n2750 N86 VDD VDD pmos w=2u l=1u
M3753 N6180 n2988 net1126 VSS nmos w=1u l=1u
M3754 net1126 n2862 VSS VSS nmos w=1u l=1u
M3755 N6180 n2988 VDD VDD pmos w=2u l=1u
M3756 N6180 n2862 VDD VDD pmos w=2u l=1u
M3757 n2988 net1127 VSS VSS nmos w=1u l=1u
M3758 net1127 n2989 VSS VSS nmos w=1u l=1u
M3759 net1127 n2990 VSS VSS nmos w=1u l=1u
M3760 net1127 n2990 net1128 VDD pmos w=2u l=1u
M3761 n2988 net1127 VDD VDD pmos w=2u l=1u
M3762 net1128 n2989 VDD VDD pmos w=2u l=1u
M3763 n2862 n2990 net1129 VSS nmos w=1u l=1u
M3764 net1129 n2989 VSS VSS nmos w=1u l=1u
M3765 n2862 n2990 VDD VDD pmos w=2u l=1u
M3766 n2862 n2989 VDD VDD pmos w=2u l=1u
M3767 n2990 n2992 net1130 VSS nmos w=1u l=1u
M3768 net1130 n2991 VSS VSS nmos w=1u l=1u
M3769 n2990 n2992 VDD VDD pmos w=2u l=1u
M3770 n2990 n2991 VDD VDD pmos w=2u l=1u
M3771 n2991 n2994 net1131 VSS nmos w=1u l=1u
M3772 net1131 n2993 VSS VSS nmos w=1u l=1u
M3773 n2991 n2994 VDD VDD pmos w=2u l=1u
M3774 n2991 n2993 VDD VDD pmos w=2u l=1u
M3775 net1132 n2864 VSS VSS nmos w=1u l=1u
M3776 net1133 n2863 VSS VSS nmos w=1u l=1u
M3777 n2989 net1134 VSS VSS nmos w=1u l=1u
M3778 net1134 n2864 net1135 VSS nmos w=1u l=1u
M3779 net1134 net1132 net1133 VSS nmos w=1u l=1u
M3780 net1135 net1133 VSS VSS nmos w=1u l=1u
M3781 net1134 net1132 net1136 VDD pmos w=2u l=1u
M3782 net1132 n2864 VDD VDD pmos w=2u l=1u
M3783 net1133 n2864 net1134 VDD pmos w=2u l=1u
M3784 net1133 n2863 VDD VDD pmos w=2u l=1u
M3785 n2989 net1134 VDD VDD pmos w=2u l=1u
M3786 net1136 net1133 VDD VDD pmos w=2u l=1u
M3787 n2864 n2996 net1137 VSS nmos w=1u l=1u
M3788 net1137 n2995 VSS VSS nmos w=1u l=1u
M3789 n2864 n2996 VDD VDD pmos w=2u l=1u
M3790 n2864 n2995 VDD VDD pmos w=2u l=1u
M3791 n2995 n2998 net1138 VSS nmos w=1u l=1u
M3792 net1138 n2997 VSS VSS nmos w=1u l=1u
M3793 n2995 n2998 VDD VDD pmos w=2u l=1u
M3794 n2995 n2997 VDD VDD pmos w=2u l=1u
M3795 net1139 n2867 VSS VSS nmos w=1u l=1u
M3796 net1140 n2868 VSS VSS nmos w=1u l=1u
M3797 n2863 net1141 VSS VSS nmos w=1u l=1u
M3798 net1141 n2867 net1142 VSS nmos w=1u l=1u
M3799 net1141 net1139 net1140 VSS nmos w=1u l=1u
M3800 net1142 net1140 VSS VSS nmos w=1u l=1u
M3801 net1141 net1139 net1143 VDD pmos w=2u l=1u
M3802 net1139 n2867 VDD VDD pmos w=2u l=1u
M3803 net1140 n2867 net1141 VDD pmos w=2u l=1u
M3804 net1140 n2868 VDD VDD pmos w=2u l=1u
M3805 n2863 net1141 VDD VDD pmos w=2u l=1u
M3806 net1143 net1140 VDD VDD pmos w=2u l=1u
M3807 n2867 net1144 VSS VSS nmos w=1u l=1u
M3808 net1145 n2866 VSS VSS nmos w=1u l=1u
M3809 net1144 n2999 net1145 VSS nmos w=1u l=1u
M3810 net1144 n2866 VDD VDD pmos w=2u l=1u
M3811 net1144 n2999 VDD VDD pmos w=2u l=1u
M3812 n2867 net1144 VDD VDD pmos w=2u l=1u
M3813 n2866 n3001 net1146 VSS nmos w=1u l=1u
M3814 net1146 n3000 VSS VSS nmos w=1u l=1u
M3815 n2866 n3001 VDD VDD pmos w=2u l=1u
M3816 n2866 n3000 VDD VDD pmos w=2u l=1u
M3817 n3001 n3003 net1147 VSS nmos w=1u l=1u
M3818 net1147 n3002 VSS VSS nmos w=1u l=1u
M3819 n3001 n3003 VDD VDD pmos w=2u l=1u
M3820 n3001 n3002 VDD VDD pmos w=2u l=1u
M3821 n3002 net1148 VSS VSS nmos w=1u l=1u
M3822 net1148 n3004 VSS VSS nmos w=1u l=1u
M3823 net1148 n3005 VSS VSS nmos w=1u l=1u
M3824 net1148 n3005 net1149 VDD pmos w=2u l=1u
M3825 n3002 net1148 VDD VDD pmos w=2u l=1u
M3826 net1149 n3004 VDD VDD pmos w=2u l=1u
M3827 net1150 n2874 VSS VSS nmos w=1u l=1u
M3828 net1151 n2875 VSS VSS nmos w=1u l=1u
M3829 n3000 net1152 VSS VSS nmos w=1u l=1u
M3830 net1152 n2874 net1153 VSS nmos w=1u l=1u
M3831 net1152 net1150 net1151 VSS nmos w=1u l=1u
M3832 net1153 net1151 VSS VSS nmos w=1u l=1u
M3833 net1152 net1150 net1154 VDD pmos w=2u l=1u
M3834 net1150 n2874 VDD VDD pmos w=2u l=1u
M3835 net1151 n2874 net1152 VDD pmos w=2u l=1u
M3836 net1151 n2875 VDD VDD pmos w=2u l=1u
M3837 n3000 net1152 VDD VDD pmos w=2u l=1u
M3838 net1154 net1151 VDD VDD pmos w=2u l=1u
M3839 n2875 n3006 VDD VDD pmos w=2u l=1u
M3840 n2875 n3006 VSS VSS nmos w=1u l=1u
M3841 n2999 n3008 net1155 VSS nmos w=1u l=1u
M3842 net1155 n3007 VSS VSS nmos w=1u l=1u
M3843 n2999 n3008 VDD VDD pmos w=2u l=1u
M3844 n2999 n3007 VDD VDD pmos w=2u l=1u
M3845 net1156 n3006 VSS VSS nmos w=1u l=1u
M3846 net1157 n2874 VSS VSS nmos w=1u l=1u
M3847 n3008 net1158 VSS VSS nmos w=1u l=1u
M3848 net1158 n3006 net1159 VSS nmos w=1u l=1u
M3849 net1158 net1156 net1157 VSS nmos w=1u l=1u
M3850 net1159 net1157 VSS VSS nmos w=1u l=1u
M3851 net1158 net1156 net1160 VDD pmos w=2u l=1u
M3852 net1156 n3006 VDD VDD pmos w=2u l=1u
M3853 net1157 n3006 net1158 VDD pmos w=2u l=1u
M3854 net1157 n2874 VDD VDD pmos w=2u l=1u
M3855 n3008 net1158 VDD VDD pmos w=2u l=1u
M3856 net1160 net1157 VDD VDD pmos w=2u l=1u
M3857 n3006 N511 net1161 VSS nmos w=1u l=1u
M3858 net1161 N86 VSS VSS nmos w=1u l=1u
M3859 n3006 N511 VDD VDD pmos w=2u l=1u
M3860 n3006 N86 VDD VDD pmos w=2u l=1u
M3861 n2874 n2873 net1162 VSS nmos w=1u l=1u
M3862 net1162 n3009 VSS VSS nmos w=1u l=1u
M3863 n2874 n2873 VDD VDD pmos w=2u l=1u
M3864 n2874 n3009 VDD VDD pmos w=2u l=1u
M3865 n2873 n3011 net1163 VSS nmos w=1u l=1u
M3866 net1163 n3010 VSS VSS nmos w=1u l=1u
M3867 n2873 n3011 VDD VDD pmos w=2u l=1u
M3868 n2873 n3010 VDD VDD pmos w=2u l=1u
M3869 n3011 n3013 net1164 VSS nmos w=1u l=1u
M3870 net1164 n3012 VSS VSS nmos w=1u l=1u
M3871 n3011 n3013 VDD VDD pmos w=2u l=1u
M3872 n3011 n3012 VDD VDD pmos w=2u l=1u
M3873 n3012 net1165 VSS VSS nmos w=1u l=1u
M3874 net1165 n3014 VSS VSS nmos w=1u l=1u
M3875 net1165 n3015 VSS VSS nmos w=1u l=1u
M3876 net1165 n3015 net1166 VDD pmos w=2u l=1u
M3877 n3012 net1165 VDD VDD pmos w=2u l=1u
M3878 net1166 n3014 VDD VDD pmos w=2u l=1u
M3879 net1167 n2884 VSS VSS nmos w=1u l=1u
M3880 net1168 n2885 VSS VSS nmos w=1u l=1u
M3881 n3010 net1169 VSS VSS nmos w=1u l=1u
M3882 net1169 n2884 net1170 VSS nmos w=1u l=1u
M3883 net1169 net1167 net1168 VSS nmos w=1u l=1u
M3884 net1170 net1168 VSS VSS nmos w=1u l=1u
M3885 net1169 net1167 net1171 VDD pmos w=2u l=1u
M3886 net1167 n2884 VDD VDD pmos w=2u l=1u
M3887 net1168 n2884 net1169 VDD pmos w=2u l=1u
M3888 net1168 n2885 VDD VDD pmos w=2u l=1u
M3889 n3010 net1169 VDD VDD pmos w=2u l=1u
M3890 net1171 net1168 VDD VDD pmos w=2u l=1u
M3891 n2885 n3016 VDD VDD pmos w=2u l=1u
M3892 n2885 n3016 VSS VSS nmos w=1u l=1u
M3893 n3009 n3018 net1172 VSS nmos w=1u l=1u
M3894 net1172 n3017 VSS VSS nmos w=1u l=1u
M3895 n3009 n3018 VDD VDD pmos w=2u l=1u
M3896 n3009 n3017 VDD VDD pmos w=2u l=1u
M3897 net1173 n3016 VSS VSS nmos w=1u l=1u
M3898 net1174 n2884 VSS VSS nmos w=1u l=1u
M3899 n3018 net1175 VSS VSS nmos w=1u l=1u
M3900 net1175 n3016 net1176 VSS nmos w=1u l=1u
M3901 net1175 net1173 net1174 VSS nmos w=1u l=1u
M3902 net1176 net1174 VSS VSS nmos w=1u l=1u
M3903 net1175 net1173 net1177 VDD pmos w=2u l=1u
M3904 net1173 n3016 VDD VDD pmos w=2u l=1u
M3905 net1174 n3016 net1175 VDD pmos w=2u l=1u
M3906 net1174 n2884 VDD VDD pmos w=2u l=1u
M3907 n3018 net1175 VDD VDD pmos w=2u l=1u
M3908 net1177 net1174 VDD VDD pmos w=2u l=1u
M3909 n3016 N494 net1178 VSS nmos w=1u l=1u
M3910 net1178 N103 VSS VSS nmos w=1u l=1u
M3911 n3016 N494 VDD VDD pmos w=2u l=1u
M3912 n3016 N103 VDD VDD pmos w=2u l=1u
M3913 n2884 n2883 net1179 VSS nmos w=1u l=1u
M3914 net1179 n3019 VSS VSS nmos w=1u l=1u
M3915 n2884 n2883 VDD VDD pmos w=2u l=1u
M3916 n2884 n3019 VDD VDD pmos w=2u l=1u
M3917 n2883 n3021 net1180 VSS nmos w=1u l=1u
M3918 net1180 n3020 VSS VSS nmos w=1u l=1u
M3919 n2883 n3021 VDD VDD pmos w=2u l=1u
M3920 n2883 n3020 VDD VDD pmos w=2u l=1u
M3921 n3021 n3023 net1181 VSS nmos w=1u l=1u
M3922 net1181 n3022 VSS VSS nmos w=1u l=1u
M3923 n3021 n3023 VDD VDD pmos w=2u l=1u
M3924 n3021 n3022 VDD VDD pmos w=2u l=1u
M3925 n3022 net1182 VSS VSS nmos w=1u l=1u
M3926 net1182 n3024 VSS VSS nmos w=1u l=1u
M3927 net1182 n3025 VSS VSS nmos w=1u l=1u
M3928 net1182 n3025 net1183 VDD pmos w=2u l=1u
M3929 n3022 net1182 VDD VDD pmos w=2u l=1u
M3930 net1183 n3024 VDD VDD pmos w=2u l=1u
M3931 net1184 n2894 VSS VSS nmos w=1u l=1u
M3932 net1185 n2895 VSS VSS nmos w=1u l=1u
M3933 n3020 net1186 VSS VSS nmos w=1u l=1u
M3934 net1186 n2894 net1187 VSS nmos w=1u l=1u
M3935 net1186 net1184 net1185 VSS nmos w=1u l=1u
M3936 net1187 net1185 VSS VSS nmos w=1u l=1u
M3937 net1186 net1184 net1188 VDD pmos w=2u l=1u
M3938 net1184 n2894 VDD VDD pmos w=2u l=1u
M3939 net1185 n2894 net1186 VDD pmos w=2u l=1u
M3940 net1185 n2895 VDD VDD pmos w=2u l=1u
M3941 n3020 net1186 VDD VDD pmos w=2u l=1u
M3942 net1188 net1185 VDD VDD pmos w=2u l=1u
M3943 n2895 n3026 VDD VDD pmos w=2u l=1u
M3944 n2895 n3026 VSS VSS nmos w=1u l=1u
M3945 n3019 n3028 net1189 VSS nmos w=1u l=1u
M3946 net1189 n3027 VSS VSS nmos w=1u l=1u
M3947 n3019 n3028 VDD VDD pmos w=2u l=1u
M3948 n3019 n3027 VDD VDD pmos w=2u l=1u
M3949 net1190 n3026 VSS VSS nmos w=1u l=1u
M3950 net1191 n2894 VSS VSS nmos w=1u l=1u
M3951 n3028 net1192 VSS VSS nmos w=1u l=1u
M3952 net1192 n3026 net1193 VSS nmos w=1u l=1u
M3953 net1192 net1190 net1191 VSS nmos w=1u l=1u
M3954 net1193 net1191 VSS VSS nmos w=1u l=1u
M3955 net1192 net1190 net1194 VDD pmos w=2u l=1u
M3956 net1190 n3026 VDD VDD pmos w=2u l=1u
M3957 net1191 n3026 net1192 VDD pmos w=2u l=1u
M3958 net1191 n2894 VDD VDD pmos w=2u l=1u
M3959 n3028 net1192 VDD VDD pmos w=2u l=1u
M3960 net1194 net1191 VDD VDD pmos w=2u l=1u
M3961 n3026 N477 net1195 VSS nmos w=1u l=1u
M3962 net1195 N120 VSS VSS nmos w=1u l=1u
M3963 n3026 N477 VDD VDD pmos w=2u l=1u
M3964 n3026 N120 VDD VDD pmos w=2u l=1u
M3965 n2894 n2893 net1196 VSS nmos w=1u l=1u
M3966 net1196 n3029 VSS VSS nmos w=1u l=1u
M3967 n2894 n2893 VDD VDD pmos w=2u l=1u
M3968 n2894 n3029 VDD VDD pmos w=2u l=1u
M3969 n2893 n3031 net1197 VSS nmos w=1u l=1u
M3970 net1197 n3030 VSS VSS nmos w=1u l=1u
M3971 n2893 n3031 VDD VDD pmos w=2u l=1u
M3972 n2893 n3030 VDD VDD pmos w=2u l=1u
M3973 n3031 n3033 net1198 VSS nmos w=1u l=1u
M3974 net1198 n3032 VSS VSS nmos w=1u l=1u
M3975 n3031 n3033 VDD VDD pmos w=2u l=1u
M3976 n3031 n3032 VDD VDD pmos w=2u l=1u
M3977 n3032 net1199 VSS VSS nmos w=1u l=1u
M3978 net1199 n3034 VSS VSS nmos w=1u l=1u
M3979 net1199 n3035 VSS VSS nmos w=1u l=1u
M3980 net1199 n3035 net1200 VDD pmos w=2u l=1u
M3981 n3032 net1199 VDD VDD pmos w=2u l=1u
M3982 net1200 n3034 VDD VDD pmos w=2u l=1u
M3983 net1201 n2904 VSS VSS nmos w=1u l=1u
M3984 net1202 n2905 VSS VSS nmos w=1u l=1u
M3985 n3030 net1203 VSS VSS nmos w=1u l=1u
M3986 net1203 n2904 net1204 VSS nmos w=1u l=1u
M3987 net1203 net1201 net1202 VSS nmos w=1u l=1u
M3988 net1204 net1202 VSS VSS nmos w=1u l=1u
M3989 net1203 net1201 net1205 VDD pmos w=2u l=1u
M3990 net1201 n2904 VDD VDD pmos w=2u l=1u
M3991 net1202 n2904 net1203 VDD pmos w=2u l=1u
M3992 net1202 n2905 VDD VDD pmos w=2u l=1u
M3993 n3030 net1203 VDD VDD pmos w=2u l=1u
M3994 net1205 net1202 VDD VDD pmos w=2u l=1u
M3995 n2905 n3036 VDD VDD pmos w=2u l=1u
M3996 n2905 n3036 VSS VSS nmos w=1u l=1u
M3997 n3029 n3038 net1206 VSS nmos w=1u l=1u
M3998 net1206 n3037 VSS VSS nmos w=1u l=1u
M3999 n3029 n3038 VDD VDD pmos w=2u l=1u
M4000 n3029 n3037 VDD VDD pmos w=2u l=1u
M4001 net1207 n3036 VSS VSS nmos w=1u l=1u
M4002 net1208 n2904 VSS VSS nmos w=1u l=1u
M4003 n3038 net1209 VSS VSS nmos w=1u l=1u
M4004 net1209 n3036 net1210 VSS nmos w=1u l=1u
M4005 net1209 net1207 net1208 VSS nmos w=1u l=1u
M4006 net1210 net1208 VSS VSS nmos w=1u l=1u
M4007 net1209 net1207 net1211 VDD pmos w=2u l=1u
M4008 net1207 n3036 VDD VDD pmos w=2u l=1u
M4009 net1208 n3036 net1209 VDD pmos w=2u l=1u
M4010 net1208 n2904 VDD VDD pmos w=2u l=1u
M4011 n3038 net1209 VDD VDD pmos w=2u l=1u
M4012 net1211 net1208 VDD VDD pmos w=2u l=1u
M4013 n3036 N460 net1212 VSS nmos w=1u l=1u
M4014 net1212 N137 VSS VSS nmos w=1u l=1u
M4015 n3036 N460 VDD VDD pmos w=2u l=1u
M4016 n3036 N137 VDD VDD pmos w=2u l=1u
M4017 n2904 n2903 net1213 VSS nmos w=1u l=1u
M4018 net1213 n3039 VSS VSS nmos w=1u l=1u
M4019 n2904 n2903 VDD VDD pmos w=2u l=1u
M4020 n2904 n3039 VDD VDD pmos w=2u l=1u
M4021 n2903 n3041 net1214 VSS nmos w=1u l=1u
M4022 net1214 n3040 VSS VSS nmos w=1u l=1u
M4023 n2903 n3041 VDD VDD pmos w=2u l=1u
M4024 n2903 n3040 VDD VDD pmos w=2u l=1u
M4025 n3041 n3043 net1215 VSS nmos w=1u l=1u
M4026 net1215 n3042 VSS VSS nmos w=1u l=1u
M4027 n3041 n3043 VDD VDD pmos w=2u l=1u
M4028 n3041 n3042 VDD VDD pmos w=2u l=1u
M4029 n3042 net1216 VSS VSS nmos w=1u l=1u
M4030 net1216 n3044 VSS VSS nmos w=1u l=1u
M4031 net1216 n3045 VSS VSS nmos w=1u l=1u
M4032 net1216 n3045 net1217 VDD pmos w=2u l=1u
M4033 n3042 net1216 VDD VDD pmos w=2u l=1u
M4034 net1217 n3044 VDD VDD pmos w=2u l=1u
M4035 net1218 n2914 VSS VSS nmos w=1u l=1u
M4036 net1219 n2915 VSS VSS nmos w=1u l=1u
M4037 n3040 net1220 VSS VSS nmos w=1u l=1u
M4038 net1220 n2914 net1221 VSS nmos w=1u l=1u
M4039 net1220 net1218 net1219 VSS nmos w=1u l=1u
M4040 net1221 net1219 VSS VSS nmos w=1u l=1u
M4041 net1220 net1218 net1222 VDD pmos w=2u l=1u
M4042 net1218 n2914 VDD VDD pmos w=2u l=1u
M4043 net1219 n2914 net1220 VDD pmos w=2u l=1u
M4044 net1219 n2915 VDD VDD pmos w=2u l=1u
M4045 n3040 net1220 VDD VDD pmos w=2u l=1u
M4046 net1222 net1219 VDD VDD pmos w=2u l=1u
M4047 n2915 n3046 VDD VDD pmos w=2u l=1u
M4048 n2915 n3046 VSS VSS nmos w=1u l=1u
M4049 n3039 n3048 net1223 VSS nmos w=1u l=1u
M4050 net1223 n3047 VSS VSS nmos w=1u l=1u
M4051 n3039 n3048 VDD VDD pmos w=2u l=1u
M4052 n3039 n3047 VDD VDD pmos w=2u l=1u
M4053 net1224 n3046 VSS VSS nmos w=1u l=1u
M4054 net1225 n2914 VSS VSS nmos w=1u l=1u
M4055 n3048 net1226 VSS VSS nmos w=1u l=1u
M4056 net1226 n3046 net1227 VSS nmos w=1u l=1u
M4057 net1226 net1224 net1225 VSS nmos w=1u l=1u
M4058 net1227 net1225 VSS VSS nmos w=1u l=1u
M4059 net1226 net1224 net1228 VDD pmos w=2u l=1u
M4060 net1224 n3046 VDD VDD pmos w=2u l=1u
M4061 net1225 n3046 net1226 VDD pmos w=2u l=1u
M4062 net1225 n2914 VDD VDD pmos w=2u l=1u
M4063 n3048 net1226 VDD VDD pmos w=2u l=1u
M4064 net1228 net1225 VDD VDD pmos w=2u l=1u
M4065 n3046 N443 net1229 VSS nmos w=1u l=1u
M4066 net1229 N154 VSS VSS nmos w=1u l=1u
M4067 n3046 N443 VDD VDD pmos w=2u l=1u
M4068 n3046 N154 VDD VDD pmos w=2u l=1u
M4069 n2914 n2913 net1230 VSS nmos w=1u l=1u
M4070 net1230 n3049 VSS VSS nmos w=1u l=1u
M4071 n2914 n2913 VDD VDD pmos w=2u l=1u
M4072 n2914 n3049 VDD VDD pmos w=2u l=1u
M4073 n2913 n3051 net1231 VSS nmos w=1u l=1u
M4074 net1231 n3050 VSS VSS nmos w=1u l=1u
M4075 n2913 n3051 VDD VDD pmos w=2u l=1u
M4076 n2913 n3050 VDD VDD pmos w=2u l=1u
M4077 n3051 n3053 net1232 VSS nmos w=1u l=1u
M4078 net1232 n3052 VSS VSS nmos w=1u l=1u
M4079 n3051 n3053 VDD VDD pmos w=2u l=1u
M4080 n3051 n3052 VDD VDD pmos w=2u l=1u
M4081 n3052 net1233 VSS VSS nmos w=1u l=1u
M4082 net1233 n3054 VSS VSS nmos w=1u l=1u
M4083 net1233 n3055 VSS VSS nmos w=1u l=1u
M4084 net1233 n3055 net1234 VDD pmos w=2u l=1u
M4085 n3052 net1233 VDD VDD pmos w=2u l=1u
M4086 net1234 n3054 VDD VDD pmos w=2u l=1u
M4087 net1235 n2924 VSS VSS nmos w=1u l=1u
M4088 net1236 n2925 VSS VSS nmos w=1u l=1u
M4089 n3050 net1237 VSS VSS nmos w=1u l=1u
M4090 net1237 n2924 net1238 VSS nmos w=1u l=1u
M4091 net1237 net1235 net1236 VSS nmos w=1u l=1u
M4092 net1238 net1236 VSS VSS nmos w=1u l=1u
M4093 net1237 net1235 net1239 VDD pmos w=2u l=1u
M4094 net1235 n2924 VDD VDD pmos w=2u l=1u
M4095 net1236 n2924 net1237 VDD pmos w=2u l=1u
M4096 net1236 n2925 VDD VDD pmos w=2u l=1u
M4097 n3050 net1237 VDD VDD pmos w=2u l=1u
M4098 net1239 net1236 VDD VDD pmos w=2u l=1u
M4099 n2925 n3056 VDD VDD pmos w=2u l=1u
M4100 n2925 n3056 VSS VSS nmos w=1u l=1u
M4101 n3049 n3058 net1240 VSS nmos w=1u l=1u
M4102 net1240 n3057 VSS VSS nmos w=1u l=1u
M4103 n3049 n3058 VDD VDD pmos w=2u l=1u
M4104 n3049 n3057 VDD VDD pmos w=2u l=1u
M4105 net1241 n3056 VSS VSS nmos w=1u l=1u
M4106 net1242 n2924 VSS VSS nmos w=1u l=1u
M4107 n3058 net1243 VSS VSS nmos w=1u l=1u
M4108 net1243 n3056 net1244 VSS nmos w=1u l=1u
M4109 net1243 net1241 net1242 VSS nmos w=1u l=1u
M4110 net1244 net1242 VSS VSS nmos w=1u l=1u
M4111 net1243 net1241 net1245 VDD pmos w=2u l=1u
M4112 net1241 n3056 VDD VDD pmos w=2u l=1u
M4113 net1242 n3056 net1243 VDD pmos w=2u l=1u
M4114 net1242 n2924 VDD VDD pmos w=2u l=1u
M4115 n3058 net1243 VDD VDD pmos w=2u l=1u
M4116 net1245 net1242 VDD VDD pmos w=2u l=1u
M4117 n3056 N426 net1246 VSS nmos w=1u l=1u
M4118 net1246 N171 VSS VSS nmos w=1u l=1u
M4119 n3056 N426 VDD VDD pmos w=2u l=1u
M4120 n3056 N171 VDD VDD pmos w=2u l=1u
M4121 n2924 n2923 net1247 VSS nmos w=1u l=1u
M4122 net1247 n3059 VSS VSS nmos w=1u l=1u
M4123 n2924 n2923 VDD VDD pmos w=2u l=1u
M4124 n2924 n3059 VDD VDD pmos w=2u l=1u
M4125 n2923 n3061 net1248 VSS nmos w=1u l=1u
M4126 net1248 n3060 VSS VSS nmos w=1u l=1u
M4127 n2923 n3061 VDD VDD pmos w=2u l=1u
M4128 n2923 n3060 VDD VDD pmos w=2u l=1u
M4129 n3061 n3063 net1249 VSS nmos w=1u l=1u
M4130 net1249 n3062 VSS VSS nmos w=1u l=1u
M4131 n3061 n3063 VDD VDD pmos w=2u l=1u
M4132 n3061 n3062 VDD VDD pmos w=2u l=1u
M4133 n3062 net1250 VSS VSS nmos w=1u l=1u
M4134 net1250 n3064 VSS VSS nmos w=1u l=1u
M4135 net1250 n3065 VSS VSS nmos w=1u l=1u
M4136 net1250 n3065 net1251 VDD pmos w=2u l=1u
M4137 n3062 net1250 VDD VDD pmos w=2u l=1u
M4138 net1251 n3064 VDD VDD pmos w=2u l=1u
M4139 net1252 n2934 VSS VSS nmos w=1u l=1u
M4140 net1253 n2935 VSS VSS nmos w=1u l=1u
M4141 n3060 net1254 VSS VSS nmos w=1u l=1u
M4142 net1254 n2934 net1255 VSS nmos w=1u l=1u
M4143 net1254 net1252 net1253 VSS nmos w=1u l=1u
M4144 net1255 net1253 VSS VSS nmos w=1u l=1u
M4145 net1254 net1252 net1256 VDD pmos w=2u l=1u
M4146 net1252 n2934 VDD VDD pmos w=2u l=1u
M4147 net1253 n2934 net1254 VDD pmos w=2u l=1u
M4148 net1253 n2935 VDD VDD pmos w=2u l=1u
M4149 n3060 net1254 VDD VDD pmos w=2u l=1u
M4150 net1256 net1253 VDD VDD pmos w=2u l=1u
M4151 n2935 n3066 VDD VDD pmos w=2u l=1u
M4152 n2935 n3066 VSS VSS nmos w=1u l=1u
M4153 n3059 n3068 net1257 VSS nmos w=1u l=1u
M4154 net1257 n3067 VSS VSS nmos w=1u l=1u
M4155 n3059 n3068 VDD VDD pmos w=2u l=1u
M4156 n3059 n3067 VDD VDD pmos w=2u l=1u
M4157 net1258 n3066 VSS VSS nmos w=1u l=1u
M4158 net1259 n2934 VSS VSS nmos w=1u l=1u
M4159 n3068 net1260 VSS VSS nmos w=1u l=1u
M4160 net1260 n3066 net1261 VSS nmos w=1u l=1u
M4161 net1260 net1258 net1259 VSS nmos w=1u l=1u
M4162 net1261 net1259 VSS VSS nmos w=1u l=1u
M4163 net1260 net1258 net1262 VDD pmos w=2u l=1u
M4164 net1258 n3066 VDD VDD pmos w=2u l=1u
M4165 net1259 n3066 net1260 VDD pmos w=2u l=1u
M4166 net1259 n2934 VDD VDD pmos w=2u l=1u
M4167 n3068 net1260 VDD VDD pmos w=2u l=1u
M4168 net1262 net1259 VDD VDD pmos w=2u l=1u
M4169 n3066 N409 net1263 VSS nmos w=1u l=1u
M4170 net1263 N188 VSS VSS nmos w=1u l=1u
M4171 n3066 N409 VDD VDD pmos w=2u l=1u
M4172 n3066 N188 VDD VDD pmos w=2u l=1u
M4173 n2934 n2933 net1264 VSS nmos w=1u l=1u
M4174 net1264 n3069 VSS VSS nmos w=1u l=1u
M4175 n2934 n2933 VDD VDD pmos w=2u l=1u
M4176 n2934 n3069 VDD VDD pmos w=2u l=1u
M4177 n2933 n3071 net1265 VSS nmos w=1u l=1u
M4178 net1265 n3070 VSS VSS nmos w=1u l=1u
M4179 n2933 n3071 VDD VDD pmos w=2u l=1u
M4180 n2933 n3070 VDD VDD pmos w=2u l=1u
M4181 n3071 n3073 net1266 VSS nmos w=1u l=1u
M4182 net1266 n3072 VSS VSS nmos w=1u l=1u
M4183 n3071 n3073 VDD VDD pmos w=2u l=1u
M4184 n3071 n3072 VDD VDD pmos w=2u l=1u
M4185 n3072 net1267 VSS VSS nmos w=1u l=1u
M4186 net1267 n3074 VSS VSS nmos w=1u l=1u
M4187 net1267 n3075 VSS VSS nmos w=1u l=1u
M4188 net1267 n3075 net1268 VDD pmos w=2u l=1u
M4189 n3072 net1267 VDD VDD pmos w=2u l=1u
M4190 net1268 n3074 VDD VDD pmos w=2u l=1u
M4191 net1269 n2944 VSS VSS nmos w=1u l=1u
M4192 net1270 n2945 VSS VSS nmos w=1u l=1u
M4193 n3070 net1271 VSS VSS nmos w=1u l=1u
M4194 net1271 n2944 net1272 VSS nmos w=1u l=1u
M4195 net1271 net1269 net1270 VSS nmos w=1u l=1u
M4196 net1272 net1270 VSS VSS nmos w=1u l=1u
M4197 net1271 net1269 net1273 VDD pmos w=2u l=1u
M4198 net1269 n2944 VDD VDD pmos w=2u l=1u
M4199 net1270 n2944 net1271 VDD pmos w=2u l=1u
M4200 net1270 n2945 VDD VDD pmos w=2u l=1u
M4201 n3070 net1271 VDD VDD pmos w=2u l=1u
M4202 net1273 net1270 VDD VDD pmos w=2u l=1u
M4203 n2944 n3076 VDD VDD pmos w=2u l=1u
M4204 n2944 n3076 VSS VSS nmos w=1u l=1u
M4205 n3069 n3078 net1274 VSS nmos w=1u l=1u
M4206 net1274 n3077 VSS VSS nmos w=1u l=1u
M4207 n3069 n3078 VDD VDD pmos w=2u l=1u
M4208 n3069 n3077 VDD VDD pmos w=2u l=1u
M4209 net1275 n2945 VSS VSS nmos w=1u l=1u
M4210 net1276 n3076 VSS VSS nmos w=1u l=1u
M4211 n3078 net1277 VSS VSS nmos w=1u l=1u
M4212 net1277 n2945 net1278 VSS nmos w=1u l=1u
M4213 net1277 net1275 net1276 VSS nmos w=1u l=1u
M4214 net1278 net1276 VSS VSS nmos w=1u l=1u
M4215 net1277 net1275 net1279 VDD pmos w=2u l=1u
M4216 net1275 n2945 VDD VDD pmos w=2u l=1u
M4217 net1276 n2945 net1277 VDD pmos w=2u l=1u
M4218 net1276 n3076 VDD VDD pmos w=2u l=1u
M4219 n3078 net1277 VDD VDD pmos w=2u l=1u
M4220 net1279 net1276 VDD VDD pmos w=2u l=1u
M4221 n2945 N392 net1280 VSS nmos w=1u l=1u
M4222 net1280 N205 VSS VSS nmos w=1u l=1u
M4223 n2945 N392 VDD VDD pmos w=2u l=1u
M4224 n2945 N205 VDD VDD pmos w=2u l=1u
M4225 n3076 n2943 net1281 VSS nmos w=1u l=1u
M4226 net1281 n3079 VSS VSS nmos w=1u l=1u
M4227 n3076 n2943 VDD VDD pmos w=2u l=1u
M4228 n3076 n3079 VDD VDD pmos w=2u l=1u
M4229 n2943 n3081 net1282 VSS nmos w=1u l=1u
M4230 net1282 n3080 VSS VSS nmos w=1u l=1u
M4231 n2943 n3081 VDD VDD pmos w=2u l=1u
M4232 n2943 n3080 VDD VDD pmos w=2u l=1u
M4233 n3081 n3083 net1283 VSS nmos w=1u l=1u
M4234 net1283 n3082 VSS VSS nmos w=1u l=1u
M4235 n3081 n3083 VDD VDD pmos w=2u l=1u
M4236 n3081 n3082 VDD VDD pmos w=2u l=1u
M4237 n3082 net1284 VSS VSS nmos w=1u l=1u
M4238 net1284 n3084 VSS VSS nmos w=1u l=1u
M4239 net1284 n3085 VSS VSS nmos w=1u l=1u
M4240 net1284 n3085 net1285 VDD pmos w=2u l=1u
M4241 n3082 net1284 VDD VDD pmos w=2u l=1u
M4242 net1285 n3084 VDD VDD pmos w=2u l=1u
M4243 net1286 n2955 VSS VSS nmos w=1u l=1u
M4244 net1287 n2956 VSS VSS nmos w=1u l=1u
M4245 n3080 net1288 VSS VSS nmos w=1u l=1u
M4246 net1288 n2955 net1289 VSS nmos w=1u l=1u
M4247 net1288 net1286 net1287 VSS nmos w=1u l=1u
M4248 net1289 net1287 VSS VSS nmos w=1u l=1u
M4249 net1288 net1286 net1290 VDD pmos w=2u l=1u
M4250 net1286 n2955 VDD VDD pmos w=2u l=1u
M4251 net1287 n2955 net1288 VDD pmos w=2u l=1u
M4252 net1287 n2956 VDD VDD pmos w=2u l=1u
M4253 n3080 net1288 VDD VDD pmos w=2u l=1u
M4254 net1290 net1287 VDD VDD pmos w=2u l=1u
M4255 n2955 n3086 VDD VDD pmos w=2u l=1u
M4256 n2955 n3086 VSS VSS nmos w=1u l=1u
M4257 n3079 n3088 net1291 VSS nmos w=1u l=1u
M4258 net1291 n3087 VSS VSS nmos w=1u l=1u
M4259 n3079 n3088 VDD VDD pmos w=2u l=1u
M4260 n3079 n3087 VDD VDD pmos w=2u l=1u
M4261 net1292 n2956 VSS VSS nmos w=1u l=1u
M4262 net1293 n3086 VSS VSS nmos w=1u l=1u
M4263 n3088 net1294 VSS VSS nmos w=1u l=1u
M4264 net1294 n2956 net1295 VSS nmos w=1u l=1u
M4265 net1294 net1292 net1293 VSS nmos w=1u l=1u
M4266 net1295 net1293 VSS VSS nmos w=1u l=1u
M4267 net1294 net1292 net1296 VDD pmos w=2u l=1u
M4268 net1292 n2956 VDD VDD pmos w=2u l=1u
M4269 net1293 n2956 net1294 VDD pmos w=2u l=1u
M4270 net1293 n3086 VDD VDD pmos w=2u l=1u
M4271 n3088 net1294 VDD VDD pmos w=2u l=1u
M4272 net1296 net1293 VDD VDD pmos w=2u l=1u
M4273 n2956 N375 net1297 VSS nmos w=1u l=1u
M4274 net1297 N222 VSS VSS nmos w=1u l=1u
M4275 n2956 N375 VDD VDD pmos w=2u l=1u
M4276 n2956 N222 VDD VDD pmos w=2u l=1u
M4277 n3086 n2953 net1298 VSS nmos w=1u l=1u
M4278 net1298 n3089 VSS VSS nmos w=1u l=1u
M4279 n3086 n2953 VDD VDD pmos w=2u l=1u
M4280 n3086 n3089 VDD VDD pmos w=2u l=1u
M4281 n2953 n3091 net1299 VSS nmos w=1u l=1u
M4282 net1299 n3090 VSS VSS nmos w=1u l=1u
M4283 n2953 n3091 VDD VDD pmos w=2u l=1u
M4284 n2953 n3090 VDD VDD pmos w=2u l=1u
M4285 n3091 n3093 net1300 VSS nmos w=1u l=1u
M4286 net1300 n3092 VSS VSS nmos w=1u l=1u
M4287 n3091 n3093 VDD VDD pmos w=2u l=1u
M4288 n3091 n3092 VDD VDD pmos w=2u l=1u
M4289 n3089 n3092 net1301 VSS nmos w=1u l=1u
M4290 net1301 n3094 VSS VSS nmos w=1u l=1u
M4291 n3089 n3092 VDD VDD pmos w=2u l=1u
M4292 n3089 n3094 VDD VDD pmos w=2u l=1u
M4293 n3092 n3096 net1302 VSS nmos w=1u l=1u
M4294 net1302 n3095 VSS VSS nmos w=1u l=1u
M4295 n3092 n3096 VDD VDD pmos w=2u l=1u
M4296 n3092 n3095 VDD VDD pmos w=2u l=1u
M4297 n3094 n3090 VSS VSS nmos w=1u l=1u
M4298 n3094 n3097 VSS VSS nmos w=1u l=1u
M4299 n3094 n3090 net1303 VDD pmos w=2u l=1u
M4300 net1303 n3097 VDD VDD pmos w=2u l=1u
M4301 n3090 net1304 VSS VSS nmos w=1u l=1u
M4302 net1305 n3098 VSS VSS nmos w=1u l=1u
M4303 net1304 n2968 net1305 VSS nmos w=1u l=1u
M4304 net1304 n3098 VDD VDD pmos w=2u l=1u
M4305 net1304 n2968 VDD VDD pmos w=2u l=1u
M4306 n3090 net1304 VDD VDD pmos w=2u l=1u
M4307 n3098 N358 net1306 VSS nmos w=1u l=1u
M4308 net1306 n3099 VSS VSS nmos w=1u l=1u
M4309 n3098 N358 VDD VDD pmos w=2u l=1u
M4310 n3098 n3099 VDD VDD pmos w=2u l=1u
M4311 n3099 n3101 VSS VSS nmos w=1u l=1u
M4312 n3099 n3100 VSS VSS nmos w=1u l=1u
M4313 n3099 n3101 net1307 VDD pmos w=2u l=1u
M4314 net1307 n3100 VDD VDD pmos w=2u l=1u
M4315 n3101 n3103 VSS VSS nmos w=1u l=1u
M4316 n3101 n3102 VSS VSS nmos w=1u l=1u
M4317 n3101 n3103 net1308 VDD pmos w=2u l=1u
M4318 net1308 n3102 VDD VDD pmos w=2u l=1u
M4319 n3103 n2270 net1309 VSS nmos w=1u l=1u
M4320 net1309 n3104 VSS VSS nmos w=1u l=1u
M4321 n3103 n2270 VDD VDD pmos w=2u l=1u
M4322 n3103 n3104 VDD VDD pmos w=2u l=1u
M4323 n3104 n3105 net1310 VSS nmos w=1u l=1u
M4324 net1310 N239 VSS VSS nmos w=1u l=1u
M4325 n3104 n3105 VDD VDD pmos w=2u l=1u
M4326 n3104 N239 VDD VDD pmos w=2u l=1u
M4327 n3102 n2971 VDD VDD pmos w=2u l=1u
M4328 n3102 n2971 VSS VSS nmos w=1u l=1u
M4329 n3100 n2971 VSS VSS nmos w=1u l=1u
M4330 n3100 N341 VSS VSS nmos w=1u l=1u
M4331 n3100 n2971 net1311 VDD pmos w=2u l=1u
M4332 net1311 N341 VDD VDD pmos w=2u l=1u
M4333 n2968 n3107 net1312 VSS nmos w=1u l=1u
M4334 net1312 n3106 VSS VSS nmos w=1u l=1u
M4335 n2968 n3107 VDD VDD pmos w=2u l=1u
M4336 n2968 n3106 VDD VDD pmos w=2u l=1u
M4337 n3107 N239 net1313 VSS nmos w=1u l=1u
M4338 net1313 N358 VSS VSS nmos w=1u l=1u
M4339 n3107 N239 VDD VDD pmos w=2u l=1u
M4340 n3107 N358 VDD VDD pmos w=2u l=1u
M4341 net1314 n2970 VSS VSS nmos w=1u l=1u
M4342 net1315 n2971 VSS VSS nmos w=1u l=1u
M4343 n3106 net1316 VSS VSS nmos w=1u l=1u
M4344 net1316 n2970 net1317 VSS nmos w=1u l=1u
M4345 net1316 net1314 net1315 VSS nmos w=1u l=1u
M4346 net1317 net1315 VSS VSS nmos w=1u l=1u
M4347 net1316 net1314 net1318 VDD pmos w=2u l=1u
M4348 net1314 n2970 VDD VDD pmos w=2u l=1u
M4349 net1315 n2970 net1316 VDD pmos w=2u l=1u
M4350 net1315 n2971 VDD VDD pmos w=2u l=1u
M4351 n3106 net1316 VDD VDD pmos w=2u l=1u
M4352 net1318 net1315 VDD VDD pmos w=2u l=1u
M4353 n2970 N256 net1319 VSS nmos w=1u l=1u
M4354 net1319 N341 VSS VSS nmos w=1u l=1u
M4355 n2970 N256 VDD VDD pmos w=2u l=1u
M4356 n2970 N341 VDD VDD pmos w=2u l=1u
M4357 n2971 n3109 net1320 VSS nmos w=1u l=1u
M4358 net1320 n3108 VSS VSS nmos w=1u l=1u
M4359 n2971 n3109 VDD VDD pmos w=2u l=1u
M4360 n2971 n3108 VDD VDD pmos w=2u l=1u
M4361 n3109 n3111 net1321 VSS nmos w=1u l=1u
M4362 net1321 n3110 VSS VSS nmos w=1u l=1u
M4363 n3109 n3111 VDD VDD pmos w=2u l=1u
M4364 n3109 n3110 VDD VDD pmos w=2u l=1u
M4365 n3097 n3093 VDD VDD pmos w=2u l=1u
M4366 n3097 n3093 VSS VSS nmos w=1u l=1u
M4367 n3087 n3113 VSS VSS nmos w=1u l=1u
M4368 n3087 n3112 VSS VSS nmos w=1u l=1u
M4369 n3087 n3113 net1322 VDD pmos w=2u l=1u
M4370 net1322 n3112 VDD VDD pmos w=2u l=1u
M4371 n3113 n3084 VSS VSS nmos w=1u l=1u
M4372 n3113 n3085 VSS VSS nmos w=1u l=1u
M4373 n3113 n3084 net1323 VDD pmos w=2u l=1u
M4374 net1323 n3085 VDD VDD pmos w=2u l=1u
M4375 n3112 n3083 VDD VDD pmos w=2u l=1u
M4376 n3112 n3083 VSS VSS nmos w=1u l=1u
M4377 n3077 n3115 VSS VSS nmos w=1u l=1u
M4378 n3077 n3114 VSS VSS nmos w=1u l=1u
M4379 n3077 n3115 net1324 VDD pmos w=2u l=1u
M4380 net1324 n3114 VDD VDD pmos w=2u l=1u
M4381 n3115 n3074 VSS VSS nmos w=1u l=1u
M4382 n3115 n3075 VSS VSS nmos w=1u l=1u
M4383 n3115 n3074 net1325 VDD pmos w=2u l=1u
M4384 net1325 n3075 VDD VDD pmos w=2u l=1u
M4385 n3114 n3073 VDD VDD pmos w=2u l=1u
M4386 n3114 n3073 VSS VSS nmos w=1u l=1u
M4387 n3067 n3117 VSS VSS nmos w=1u l=1u
M4388 n3067 n3116 VSS VSS nmos w=1u l=1u
M4389 n3067 n3117 net1326 VDD pmos w=2u l=1u
M4390 net1326 n3116 VDD VDD pmos w=2u l=1u
M4391 n3117 n3064 VSS VSS nmos w=1u l=1u
M4392 n3117 n3065 VSS VSS nmos w=1u l=1u
M4393 n3117 n3064 net1327 VDD pmos w=2u l=1u
M4394 net1327 n3065 VDD VDD pmos w=2u l=1u
M4395 n3116 n3063 VDD VDD pmos w=2u l=1u
M4396 n3116 n3063 VSS VSS nmos w=1u l=1u
M4397 n3057 n3119 VSS VSS nmos w=1u l=1u
M4398 n3057 n3118 VSS VSS nmos w=1u l=1u
M4399 n3057 n3119 net1328 VDD pmos w=2u l=1u
M4400 net1328 n3118 VDD VDD pmos w=2u l=1u
M4401 n3119 n3054 VSS VSS nmos w=1u l=1u
M4402 n3119 n3055 VSS VSS nmos w=1u l=1u
M4403 n3119 n3054 net1329 VDD pmos w=2u l=1u
M4404 net1329 n3055 VDD VDD pmos w=2u l=1u
M4405 n3118 n3053 VDD VDD pmos w=2u l=1u
M4406 n3118 n3053 VSS VSS nmos w=1u l=1u
M4407 n3047 n3121 VSS VSS nmos w=1u l=1u
M4408 n3047 n3120 VSS VSS nmos w=1u l=1u
M4409 n3047 n3121 net1330 VDD pmos w=2u l=1u
M4410 net1330 n3120 VDD VDD pmos w=2u l=1u
M4411 n3121 n3044 VSS VSS nmos w=1u l=1u
M4412 n3121 n3045 VSS VSS nmos w=1u l=1u
M4413 n3121 n3044 net1331 VDD pmos w=2u l=1u
M4414 net1331 n3045 VDD VDD pmos w=2u l=1u
M4415 n3120 n3043 VDD VDD pmos w=2u l=1u
M4416 n3120 n3043 VSS VSS nmos w=1u l=1u
M4417 n3037 n3123 VSS VSS nmos w=1u l=1u
M4418 n3037 n3122 VSS VSS nmos w=1u l=1u
M4419 n3037 n3123 net1332 VDD pmos w=2u l=1u
M4420 net1332 n3122 VDD VDD pmos w=2u l=1u
M4421 n3123 n3034 VSS VSS nmos w=1u l=1u
M4422 n3123 n3035 VSS VSS nmos w=1u l=1u
M4423 n3123 n3034 net1333 VDD pmos w=2u l=1u
M4424 net1333 n3035 VDD VDD pmos w=2u l=1u
M4425 n3122 n3033 VDD VDD pmos w=2u l=1u
M4426 n3122 n3033 VSS VSS nmos w=1u l=1u
M4427 n3027 n3125 VSS VSS nmos w=1u l=1u
M4428 n3027 n3124 VSS VSS nmos w=1u l=1u
M4429 n3027 n3125 net1334 VDD pmos w=2u l=1u
M4430 net1334 n3124 VDD VDD pmos w=2u l=1u
M4431 n3125 n3024 VSS VSS nmos w=1u l=1u
M4432 n3125 n3025 VSS VSS nmos w=1u l=1u
M4433 n3125 n3024 net1335 VDD pmos w=2u l=1u
M4434 net1335 n3025 VDD VDD pmos w=2u l=1u
M4435 n3124 n3023 VDD VDD pmos w=2u l=1u
M4436 n3124 n3023 VSS VSS nmos w=1u l=1u
M4437 n3017 n3127 VSS VSS nmos w=1u l=1u
M4438 n3017 n3126 VSS VSS nmos w=1u l=1u
M4439 n3017 n3127 net1336 VDD pmos w=2u l=1u
M4440 net1336 n3126 VDD VDD pmos w=2u l=1u
M4441 n3127 n3014 VSS VSS nmos w=1u l=1u
M4442 n3127 n3015 VSS VSS nmos w=1u l=1u
M4443 n3127 n3014 net1337 VDD pmos w=2u l=1u
M4444 net1337 n3015 VDD VDD pmos w=2u l=1u
M4445 n3126 n3013 VDD VDD pmos w=2u l=1u
M4446 n3126 n3013 VSS VSS nmos w=1u l=1u
M4447 n3007 n3129 VSS VSS nmos w=1u l=1u
M4448 n3007 n3128 VSS VSS nmos w=1u l=1u
M4449 n3007 n3129 net1338 VDD pmos w=2u l=1u
M4450 net1338 n3128 VDD VDD pmos w=2u l=1u
M4451 n3129 n3004 VSS VSS nmos w=1u l=1u
M4452 n3129 n3005 VSS VSS nmos w=1u l=1u
M4453 n3129 n3004 net1339 VDD pmos w=2u l=1u
M4454 net1339 n3005 VDD VDD pmos w=2u l=1u
M4455 n3128 n3003 VDD VDD pmos w=2u l=1u
M4456 n3128 n3003 VSS VSS nmos w=1u l=1u
M4457 n2868 N528 net1340 VSS nmos w=1u l=1u
M4458 net1340 N69 VSS VSS nmos w=1u l=1u
M4459 n2868 N528 VDD VDD pmos w=2u l=1u
M4460 n2868 N69 VDD VDD pmos w=2u l=1u
M4461 N6170 n3130 net1341 VSS nmos w=1u l=1u
M4462 net1341 n2992 VSS VSS nmos w=1u l=1u
M4463 N6170 n3130 VDD VDD pmos w=2u l=1u
M4464 N6170 n2992 VDD VDD pmos w=2u l=1u
M4465 n3130 net1342 VSS VSS nmos w=1u l=1u
M4466 net1342 n3131 VSS VSS nmos w=1u l=1u
M4467 net1342 n3132 VSS VSS nmos w=1u l=1u
M4468 net1342 n3132 net1343 VDD pmos w=2u l=1u
M4469 n3130 net1342 VDD VDD pmos w=2u l=1u
M4470 net1343 n3131 VDD VDD pmos w=2u l=1u
M4471 n2992 n3132 net1344 VSS nmos w=1u l=1u
M4472 net1344 n3131 VSS VSS nmos w=1u l=1u
M4473 n2992 n3132 VDD VDD pmos w=2u l=1u
M4474 n2992 n3131 VDD VDD pmos w=2u l=1u
M4475 n3132 n3134 net1345 VSS nmos w=1u l=1u
M4476 net1345 n3133 VSS VSS nmos w=1u l=1u
M4477 n3132 n3134 VDD VDD pmos w=2u l=1u
M4478 n3132 n3133 VDD VDD pmos w=2u l=1u
M4479 n3133 n3136 net1346 VSS nmos w=1u l=1u
M4480 net1346 n3135 VSS VSS nmos w=1u l=1u
M4481 n3133 n3136 VDD VDD pmos w=2u l=1u
M4482 n3133 n3135 VDD VDD pmos w=2u l=1u
M4483 net1347 n2994 VSS VSS nmos w=1u l=1u
M4484 net1348 n2993 VSS VSS nmos w=1u l=1u
M4485 n3131 net1349 VSS VSS nmos w=1u l=1u
M4486 net1349 n2994 net1350 VSS nmos w=1u l=1u
M4487 net1349 net1347 net1348 VSS nmos w=1u l=1u
M4488 net1350 net1348 VSS VSS nmos w=1u l=1u
M4489 net1349 net1347 net1351 VDD pmos w=2u l=1u
M4490 net1347 n2994 VDD VDD pmos w=2u l=1u
M4491 net1348 n2994 net1349 VDD pmos w=2u l=1u
M4492 net1348 n2993 VDD VDD pmos w=2u l=1u
M4493 n3131 net1349 VDD VDD pmos w=2u l=1u
M4494 net1351 net1348 VDD VDD pmos w=2u l=1u
M4495 n2994 n3138 net1352 VSS nmos w=1u l=1u
M4496 net1352 n3137 VSS VSS nmos w=1u l=1u
M4497 n2994 n3138 VDD VDD pmos w=2u l=1u
M4498 n2994 n3137 VDD VDD pmos w=2u l=1u
M4499 n3137 n3140 net1353 VSS nmos w=1u l=1u
M4500 net1353 n3139 VSS VSS nmos w=1u l=1u
M4501 n3137 n3140 VDD VDD pmos w=2u l=1u
M4502 n3137 n3139 VDD VDD pmos w=2u l=1u
M4503 net1354 n2997 VSS VSS nmos w=1u l=1u
M4504 net1355 n2998 VSS VSS nmos w=1u l=1u
M4505 n2993 net1356 VSS VSS nmos w=1u l=1u
M4506 net1356 n2997 net1357 VSS nmos w=1u l=1u
M4507 net1356 net1354 net1355 VSS nmos w=1u l=1u
M4508 net1357 net1355 VSS VSS nmos w=1u l=1u
M4509 net1356 net1354 net1358 VDD pmos w=2u l=1u
M4510 net1354 n2997 VDD VDD pmos w=2u l=1u
M4511 net1355 n2997 net1356 VDD pmos w=2u l=1u
M4512 net1355 n2998 VDD VDD pmos w=2u l=1u
M4513 n2993 net1356 VDD VDD pmos w=2u l=1u
M4514 net1358 net1355 VDD VDD pmos w=2u l=1u
M4515 n2997 net1359 VSS VSS nmos w=1u l=1u
M4516 net1360 n2996 VSS VSS nmos w=1u l=1u
M4517 net1359 n3141 net1360 VSS nmos w=1u l=1u
M4518 net1359 n2996 VDD VDD pmos w=2u l=1u
M4519 net1359 n3141 VDD VDD pmos w=2u l=1u
M4520 n2997 net1359 VDD VDD pmos w=2u l=1u
M4521 n2996 n3143 net1361 VSS nmos w=1u l=1u
M4522 net1361 n3142 VSS VSS nmos w=1u l=1u
M4523 n2996 n3143 VDD VDD pmos w=2u l=1u
M4524 n2996 n3142 VDD VDD pmos w=2u l=1u
M4525 n3143 n3145 net1362 VSS nmos w=1u l=1u
M4526 net1362 n3144 VSS VSS nmos w=1u l=1u
M4527 n3143 n3145 VDD VDD pmos w=2u l=1u
M4528 n3143 n3144 VDD VDD pmos w=2u l=1u
M4529 n3144 net1363 VSS VSS nmos w=1u l=1u
M4530 net1363 n3146 VSS VSS nmos w=1u l=1u
M4531 net1363 n3147 VSS VSS nmos w=1u l=1u
M4532 net1363 n3147 net1364 VDD pmos w=2u l=1u
M4533 n3144 net1363 VDD VDD pmos w=2u l=1u
M4534 net1364 n3146 VDD VDD pmos w=2u l=1u
M4535 net1365 n3004 VSS VSS nmos w=1u l=1u
M4536 net1366 n3005 VSS VSS nmos w=1u l=1u
M4537 n3142 net1367 VSS VSS nmos w=1u l=1u
M4538 net1367 n3004 net1368 VSS nmos w=1u l=1u
M4539 net1367 net1365 net1366 VSS nmos w=1u l=1u
M4540 net1368 net1366 VSS VSS nmos w=1u l=1u
M4541 net1367 net1365 net1369 VDD pmos w=2u l=1u
M4542 net1365 n3004 VDD VDD pmos w=2u l=1u
M4543 net1366 n3004 net1367 VDD pmos w=2u l=1u
M4544 net1366 n3005 VDD VDD pmos w=2u l=1u
M4545 n3142 net1367 VDD VDD pmos w=2u l=1u
M4546 net1369 net1366 VDD VDD pmos w=2u l=1u
M4547 n3005 n3148 VDD VDD pmos w=2u l=1u
M4548 n3005 n3148 VSS VSS nmos w=1u l=1u
M4549 n3141 n3150 net1370 VSS nmos w=1u l=1u
M4550 net1370 n3149 VSS VSS nmos w=1u l=1u
M4551 n3141 n3150 VDD VDD pmos w=2u l=1u
M4552 n3141 n3149 VDD VDD pmos w=2u l=1u
M4553 net1371 n3148 VSS VSS nmos w=1u l=1u
M4554 net1372 n3004 VSS VSS nmos w=1u l=1u
M4555 n3150 net1373 VSS VSS nmos w=1u l=1u
M4556 net1373 n3148 net1374 VSS nmos w=1u l=1u
M4557 net1373 net1371 net1372 VSS nmos w=1u l=1u
M4558 net1374 net1372 VSS VSS nmos w=1u l=1u
M4559 net1373 net1371 net1375 VDD pmos w=2u l=1u
M4560 net1371 n3148 VDD VDD pmos w=2u l=1u
M4561 net1372 n3148 net1373 VDD pmos w=2u l=1u
M4562 net1372 n3004 VDD VDD pmos w=2u l=1u
M4563 n3150 net1373 VDD VDD pmos w=2u l=1u
M4564 net1375 net1372 VDD VDD pmos w=2u l=1u
M4565 n3148 N511 net1376 VSS nmos w=1u l=1u
M4566 net1376 N69 VSS VSS nmos w=1u l=1u
M4567 n3148 N511 VDD VDD pmos w=2u l=1u
M4568 n3148 N69 VDD VDD pmos w=2u l=1u
M4569 n3004 n3003 net1377 VSS nmos w=1u l=1u
M4570 net1377 n3151 VSS VSS nmos w=1u l=1u
M4571 n3004 n3003 VDD VDD pmos w=2u l=1u
M4572 n3004 n3151 VDD VDD pmos w=2u l=1u
M4573 n3003 n3153 net1378 VSS nmos w=1u l=1u
M4574 net1378 n3152 VSS VSS nmos w=1u l=1u
M4575 n3003 n3153 VDD VDD pmos w=2u l=1u
M4576 n3003 n3152 VDD VDD pmos w=2u l=1u
M4577 n3153 n3155 net1379 VSS nmos w=1u l=1u
M4578 net1379 n3154 VSS VSS nmos w=1u l=1u
M4579 n3153 n3155 VDD VDD pmos w=2u l=1u
M4580 n3153 n3154 VDD VDD pmos w=2u l=1u
M4581 n3154 net1380 VSS VSS nmos w=1u l=1u
M4582 net1380 n3156 VSS VSS nmos w=1u l=1u
M4583 net1380 n3157 VSS VSS nmos w=1u l=1u
M4584 net1380 n3157 net1381 VDD pmos w=2u l=1u
M4585 n3154 net1380 VDD VDD pmos w=2u l=1u
M4586 net1381 n3156 VDD VDD pmos w=2u l=1u
M4587 net1382 n3014 VSS VSS nmos w=1u l=1u
M4588 net1383 n3015 VSS VSS nmos w=1u l=1u
M4589 n3152 net1384 VSS VSS nmos w=1u l=1u
M4590 net1384 n3014 net1385 VSS nmos w=1u l=1u
M4591 net1384 net1382 net1383 VSS nmos w=1u l=1u
M4592 net1385 net1383 VSS VSS nmos w=1u l=1u
M4593 net1384 net1382 net1386 VDD pmos w=2u l=1u
M4594 net1382 n3014 VDD VDD pmos w=2u l=1u
M4595 net1383 n3014 net1384 VDD pmos w=2u l=1u
M4596 net1383 n3015 VDD VDD pmos w=2u l=1u
M4597 n3152 net1384 VDD VDD pmos w=2u l=1u
M4598 net1386 net1383 VDD VDD pmos w=2u l=1u
M4599 n3015 n3158 VDD VDD pmos w=2u l=1u
M4600 n3015 n3158 VSS VSS nmos w=1u l=1u
M4601 n3151 n3160 net1387 VSS nmos w=1u l=1u
M4602 net1387 n3159 VSS VSS nmos w=1u l=1u
M4603 n3151 n3160 VDD VDD pmos w=2u l=1u
M4604 n3151 n3159 VDD VDD pmos w=2u l=1u
M4605 net1388 n3158 VSS VSS nmos w=1u l=1u
M4606 net1389 n3014 VSS VSS nmos w=1u l=1u
M4607 n3160 net1390 VSS VSS nmos w=1u l=1u
M4608 net1390 n3158 net1391 VSS nmos w=1u l=1u
M4609 net1390 net1388 net1389 VSS nmos w=1u l=1u
M4610 net1391 net1389 VSS VSS nmos w=1u l=1u
M4611 net1390 net1388 net1392 VDD pmos w=2u l=1u
M4612 net1388 n3158 VDD VDD pmos w=2u l=1u
M4613 net1389 n3158 net1390 VDD pmos w=2u l=1u
M4614 net1389 n3014 VDD VDD pmos w=2u l=1u
M4615 n3160 net1390 VDD VDD pmos w=2u l=1u
M4616 net1392 net1389 VDD VDD pmos w=2u l=1u
M4617 n3158 N494 net1393 VSS nmos w=1u l=1u
M4618 net1393 N86 VSS VSS nmos w=1u l=1u
M4619 n3158 N494 VDD VDD pmos w=2u l=1u
M4620 n3158 N86 VDD VDD pmos w=2u l=1u
M4621 n3014 n3013 net1394 VSS nmos w=1u l=1u
M4622 net1394 n3161 VSS VSS nmos w=1u l=1u
M4623 n3014 n3013 VDD VDD pmos w=2u l=1u
M4624 n3014 n3161 VDD VDD pmos w=2u l=1u
M4625 n3013 n3163 net1395 VSS nmos w=1u l=1u
M4626 net1395 n3162 VSS VSS nmos w=1u l=1u
M4627 n3013 n3163 VDD VDD pmos w=2u l=1u
M4628 n3013 n3162 VDD VDD pmos w=2u l=1u
M4629 n3163 n3165 net1396 VSS nmos w=1u l=1u
M4630 net1396 n3164 VSS VSS nmos w=1u l=1u
M4631 n3163 n3165 VDD VDD pmos w=2u l=1u
M4632 n3163 n3164 VDD VDD pmos w=2u l=1u
M4633 n3164 net1397 VSS VSS nmos w=1u l=1u
M4634 net1397 n3166 VSS VSS nmos w=1u l=1u
M4635 net1397 n3167 VSS VSS nmos w=1u l=1u
M4636 net1397 n3167 net1398 VDD pmos w=2u l=1u
M4637 n3164 net1397 VDD VDD pmos w=2u l=1u
M4638 net1398 n3166 VDD VDD pmos w=2u l=1u
M4639 net1399 n3024 VSS VSS nmos w=1u l=1u
M4640 net1400 n3025 VSS VSS nmos w=1u l=1u
M4641 n3162 net1401 VSS VSS nmos w=1u l=1u
M4642 net1401 n3024 net1402 VSS nmos w=1u l=1u
M4643 net1401 net1399 net1400 VSS nmos w=1u l=1u
M4644 net1402 net1400 VSS VSS nmos w=1u l=1u
M4645 net1401 net1399 net1403 VDD pmos w=2u l=1u
M4646 net1399 n3024 VDD VDD pmos w=2u l=1u
M4647 net1400 n3024 net1401 VDD pmos w=2u l=1u
M4648 net1400 n3025 VDD VDD pmos w=2u l=1u
M4649 n3162 net1401 VDD VDD pmos w=2u l=1u
M4650 net1403 net1400 VDD VDD pmos w=2u l=1u
M4651 n3025 n3168 VDD VDD pmos w=2u l=1u
M4652 n3025 n3168 VSS VSS nmos w=1u l=1u
M4653 n3161 n3170 net1404 VSS nmos w=1u l=1u
M4654 net1404 n3169 VSS VSS nmos w=1u l=1u
M4655 n3161 n3170 VDD VDD pmos w=2u l=1u
M4656 n3161 n3169 VDD VDD pmos w=2u l=1u
M4657 net1405 n3168 VSS VSS nmos w=1u l=1u
M4658 net1406 n3024 VSS VSS nmos w=1u l=1u
M4659 n3170 net1407 VSS VSS nmos w=1u l=1u
M4660 net1407 n3168 net1408 VSS nmos w=1u l=1u
M4661 net1407 net1405 net1406 VSS nmos w=1u l=1u
M4662 net1408 net1406 VSS VSS nmos w=1u l=1u
M4663 net1407 net1405 net1409 VDD pmos w=2u l=1u
M4664 net1405 n3168 VDD VDD pmos w=2u l=1u
M4665 net1406 n3168 net1407 VDD pmos w=2u l=1u
M4666 net1406 n3024 VDD VDD pmos w=2u l=1u
M4667 n3170 net1407 VDD VDD pmos w=2u l=1u
M4668 net1409 net1406 VDD VDD pmos w=2u l=1u
M4669 n3168 N477 net1410 VSS nmos w=1u l=1u
M4670 net1410 N103 VSS VSS nmos w=1u l=1u
M4671 n3168 N477 VDD VDD pmos w=2u l=1u
M4672 n3168 N103 VDD VDD pmos w=2u l=1u
M4673 n3024 n3023 net1411 VSS nmos w=1u l=1u
M4674 net1411 n3171 VSS VSS nmos w=1u l=1u
M4675 n3024 n3023 VDD VDD pmos w=2u l=1u
M4676 n3024 n3171 VDD VDD pmos w=2u l=1u
M4677 n3023 n3173 net1412 VSS nmos w=1u l=1u
M4678 net1412 n3172 VSS VSS nmos w=1u l=1u
M4679 n3023 n3173 VDD VDD pmos w=2u l=1u
M4680 n3023 n3172 VDD VDD pmos w=2u l=1u
M4681 n3173 n3175 net1413 VSS nmos w=1u l=1u
M4682 net1413 n3174 VSS VSS nmos w=1u l=1u
M4683 n3173 n3175 VDD VDD pmos w=2u l=1u
M4684 n3173 n3174 VDD VDD pmos w=2u l=1u
M4685 n3174 net1414 VSS VSS nmos w=1u l=1u
M4686 net1414 n3176 VSS VSS nmos w=1u l=1u
M4687 net1414 n3177 VSS VSS nmos w=1u l=1u
M4688 net1414 n3177 net1415 VDD pmos w=2u l=1u
M4689 n3174 net1414 VDD VDD pmos w=2u l=1u
M4690 net1415 n3176 VDD VDD pmos w=2u l=1u
M4691 net1416 n3034 VSS VSS nmos w=1u l=1u
M4692 net1417 n3035 VSS VSS nmos w=1u l=1u
M4693 n3172 net1418 VSS VSS nmos w=1u l=1u
M4694 net1418 n3034 net1419 VSS nmos w=1u l=1u
M4695 net1418 net1416 net1417 VSS nmos w=1u l=1u
M4696 net1419 net1417 VSS VSS nmos w=1u l=1u
M4697 net1418 net1416 net1420 VDD pmos w=2u l=1u
M4698 net1416 n3034 VDD VDD pmos w=2u l=1u
M4699 net1417 n3034 net1418 VDD pmos w=2u l=1u
M4700 net1417 n3035 VDD VDD pmos w=2u l=1u
M4701 n3172 net1418 VDD VDD pmos w=2u l=1u
M4702 net1420 net1417 VDD VDD pmos w=2u l=1u
M4703 n3035 n3178 VDD VDD pmos w=2u l=1u
M4704 n3035 n3178 VSS VSS nmos w=1u l=1u
M4705 n3171 n3180 net1421 VSS nmos w=1u l=1u
M4706 net1421 n3179 VSS VSS nmos w=1u l=1u
M4707 n3171 n3180 VDD VDD pmos w=2u l=1u
M4708 n3171 n3179 VDD VDD pmos w=2u l=1u
M4709 net1422 n3178 VSS VSS nmos w=1u l=1u
M4710 net1423 n3034 VSS VSS nmos w=1u l=1u
M4711 n3180 net1424 VSS VSS nmos w=1u l=1u
M4712 net1424 n3178 net1425 VSS nmos w=1u l=1u
M4713 net1424 net1422 net1423 VSS nmos w=1u l=1u
M4714 net1425 net1423 VSS VSS nmos w=1u l=1u
M4715 net1424 net1422 net1426 VDD pmos w=2u l=1u
M4716 net1422 n3178 VDD VDD pmos w=2u l=1u
M4717 net1423 n3178 net1424 VDD pmos w=2u l=1u
M4718 net1423 n3034 VDD VDD pmos w=2u l=1u
M4719 n3180 net1424 VDD VDD pmos w=2u l=1u
M4720 net1426 net1423 VDD VDD pmos w=2u l=1u
M4721 n3178 N460 net1427 VSS nmos w=1u l=1u
M4722 net1427 N120 VSS VSS nmos w=1u l=1u
M4723 n3178 N460 VDD VDD pmos w=2u l=1u
M4724 n3178 N120 VDD VDD pmos w=2u l=1u
M4725 n3034 n3033 net1428 VSS nmos w=1u l=1u
M4726 net1428 n3181 VSS VSS nmos w=1u l=1u
M4727 n3034 n3033 VDD VDD pmos w=2u l=1u
M4728 n3034 n3181 VDD VDD pmos w=2u l=1u
M4729 n3033 n3183 net1429 VSS nmos w=1u l=1u
M4730 net1429 n3182 VSS VSS nmos w=1u l=1u
M4731 n3033 n3183 VDD VDD pmos w=2u l=1u
M4732 n3033 n3182 VDD VDD pmos w=2u l=1u
M4733 n3183 n3185 net1430 VSS nmos w=1u l=1u
M4734 net1430 n3184 VSS VSS nmos w=1u l=1u
M4735 n3183 n3185 VDD VDD pmos w=2u l=1u
M4736 n3183 n3184 VDD VDD pmos w=2u l=1u
M4737 n3184 net1431 VSS VSS nmos w=1u l=1u
M4738 net1431 n3186 VSS VSS nmos w=1u l=1u
M4739 net1431 n3187 VSS VSS nmos w=1u l=1u
M4740 net1431 n3187 net1432 VDD pmos w=2u l=1u
M4741 n3184 net1431 VDD VDD pmos w=2u l=1u
M4742 net1432 n3186 VDD VDD pmos w=2u l=1u
M4743 net1433 n3044 VSS VSS nmos w=1u l=1u
M4744 net1434 n3045 VSS VSS nmos w=1u l=1u
M4745 n3182 net1435 VSS VSS nmos w=1u l=1u
M4746 net1435 n3044 net1436 VSS nmos w=1u l=1u
M4747 net1435 net1433 net1434 VSS nmos w=1u l=1u
M4748 net1436 net1434 VSS VSS nmos w=1u l=1u
M4749 net1435 net1433 net1437 VDD pmos w=2u l=1u
M4750 net1433 n3044 VDD VDD pmos w=2u l=1u
M4751 net1434 n3044 net1435 VDD pmos w=2u l=1u
M4752 net1434 n3045 VDD VDD pmos w=2u l=1u
M4753 n3182 net1435 VDD VDD pmos w=2u l=1u
M4754 net1437 net1434 VDD VDD pmos w=2u l=1u
M4755 n3045 n3188 VDD VDD pmos w=2u l=1u
M4756 n3045 n3188 VSS VSS nmos w=1u l=1u
M4757 n3181 n3190 net1438 VSS nmos w=1u l=1u
M4758 net1438 n3189 VSS VSS nmos w=1u l=1u
M4759 n3181 n3190 VDD VDD pmos w=2u l=1u
M4760 n3181 n3189 VDD VDD pmos w=2u l=1u
M4761 net1439 n3188 VSS VSS nmos w=1u l=1u
M4762 net1440 n3044 VSS VSS nmos w=1u l=1u
M4763 n3190 net1441 VSS VSS nmos w=1u l=1u
M4764 net1441 n3188 net1442 VSS nmos w=1u l=1u
M4765 net1441 net1439 net1440 VSS nmos w=1u l=1u
M4766 net1442 net1440 VSS VSS nmos w=1u l=1u
M4767 net1441 net1439 net1443 VDD pmos w=2u l=1u
M4768 net1439 n3188 VDD VDD pmos w=2u l=1u
M4769 net1440 n3188 net1441 VDD pmos w=2u l=1u
M4770 net1440 n3044 VDD VDD pmos w=2u l=1u
M4771 n3190 net1441 VDD VDD pmos w=2u l=1u
M4772 net1443 net1440 VDD VDD pmos w=2u l=1u
M4773 n3188 N443 net1444 VSS nmos w=1u l=1u
M4774 net1444 N137 VSS VSS nmos w=1u l=1u
M4775 n3188 N443 VDD VDD pmos w=2u l=1u
M4776 n3188 N137 VDD VDD pmos w=2u l=1u
M4777 n3044 n3043 net1445 VSS nmos w=1u l=1u
M4778 net1445 n3191 VSS VSS nmos w=1u l=1u
M4779 n3044 n3043 VDD VDD pmos w=2u l=1u
M4780 n3044 n3191 VDD VDD pmos w=2u l=1u
M4781 n3043 n3193 net1446 VSS nmos w=1u l=1u
M4782 net1446 n3192 VSS VSS nmos w=1u l=1u
M4783 n3043 n3193 VDD VDD pmos w=2u l=1u
M4784 n3043 n3192 VDD VDD pmos w=2u l=1u
M4785 n3193 n3195 net1447 VSS nmos w=1u l=1u
M4786 net1447 n3194 VSS VSS nmos w=1u l=1u
M4787 n3193 n3195 VDD VDD pmos w=2u l=1u
M4788 n3193 n3194 VDD VDD pmos w=2u l=1u
M4789 n3194 net1448 VSS VSS nmos w=1u l=1u
M4790 net1448 n3196 VSS VSS nmos w=1u l=1u
M4791 net1448 n3197 VSS VSS nmos w=1u l=1u
M4792 net1448 n3197 net1449 VDD pmos w=2u l=1u
M4793 n3194 net1448 VDD VDD pmos w=2u l=1u
M4794 net1449 n3196 VDD VDD pmos w=2u l=1u
M4795 net1450 n3054 VSS VSS nmos w=1u l=1u
M4796 net1451 n3055 VSS VSS nmos w=1u l=1u
M4797 n3192 net1452 VSS VSS nmos w=1u l=1u
M4798 net1452 n3054 net1453 VSS nmos w=1u l=1u
M4799 net1452 net1450 net1451 VSS nmos w=1u l=1u
M4800 net1453 net1451 VSS VSS nmos w=1u l=1u
M4801 net1452 net1450 net1454 VDD pmos w=2u l=1u
M4802 net1450 n3054 VDD VDD pmos w=2u l=1u
M4803 net1451 n3054 net1452 VDD pmos w=2u l=1u
M4804 net1451 n3055 VDD VDD pmos w=2u l=1u
M4805 n3192 net1452 VDD VDD pmos w=2u l=1u
M4806 net1454 net1451 VDD VDD pmos w=2u l=1u
M4807 n3055 n3198 VDD VDD pmos w=2u l=1u
M4808 n3055 n3198 VSS VSS nmos w=1u l=1u
M4809 n3191 n3200 net1455 VSS nmos w=1u l=1u
M4810 net1455 n3199 VSS VSS nmos w=1u l=1u
M4811 n3191 n3200 VDD VDD pmos w=2u l=1u
M4812 n3191 n3199 VDD VDD pmos w=2u l=1u
M4813 net1456 n3198 VSS VSS nmos w=1u l=1u
M4814 net1457 n3054 VSS VSS nmos w=1u l=1u
M4815 n3200 net1458 VSS VSS nmos w=1u l=1u
M4816 net1458 n3198 net1459 VSS nmos w=1u l=1u
M4817 net1458 net1456 net1457 VSS nmos w=1u l=1u
M4818 net1459 net1457 VSS VSS nmos w=1u l=1u
M4819 net1458 net1456 net1460 VDD pmos w=2u l=1u
M4820 net1456 n3198 VDD VDD pmos w=2u l=1u
M4821 net1457 n3198 net1458 VDD pmos w=2u l=1u
M4822 net1457 n3054 VDD VDD pmos w=2u l=1u
M4823 n3200 net1458 VDD VDD pmos w=2u l=1u
M4824 net1460 net1457 VDD VDD pmos w=2u l=1u
M4825 n3198 N426 net1461 VSS nmos w=1u l=1u
M4826 net1461 N154 VSS VSS nmos w=1u l=1u
M4827 n3198 N426 VDD VDD pmos w=2u l=1u
M4828 n3198 N154 VDD VDD pmos w=2u l=1u
M4829 n3054 n3053 net1462 VSS nmos w=1u l=1u
M4830 net1462 n3201 VSS VSS nmos w=1u l=1u
M4831 n3054 n3053 VDD VDD pmos w=2u l=1u
M4832 n3054 n3201 VDD VDD pmos w=2u l=1u
M4833 n3053 n3203 net1463 VSS nmos w=1u l=1u
M4834 net1463 n3202 VSS VSS nmos w=1u l=1u
M4835 n3053 n3203 VDD VDD pmos w=2u l=1u
M4836 n3053 n3202 VDD VDD pmos w=2u l=1u
M4837 n3203 n3205 net1464 VSS nmos w=1u l=1u
M4838 net1464 n3204 VSS VSS nmos w=1u l=1u
M4839 n3203 n3205 VDD VDD pmos w=2u l=1u
M4840 n3203 n3204 VDD VDD pmos w=2u l=1u
M4841 n3204 net1465 VSS VSS nmos w=1u l=1u
M4842 net1465 n3206 VSS VSS nmos w=1u l=1u
M4843 net1465 n3207 VSS VSS nmos w=1u l=1u
M4844 net1465 n3207 net1466 VDD pmos w=2u l=1u
M4845 n3204 net1465 VDD VDD pmos w=2u l=1u
M4846 net1466 n3206 VDD VDD pmos w=2u l=1u
M4847 net1467 n3064 VSS VSS nmos w=1u l=1u
M4848 net1468 n3065 VSS VSS nmos w=1u l=1u
M4849 n3202 net1469 VSS VSS nmos w=1u l=1u
M4850 net1469 n3064 net1470 VSS nmos w=1u l=1u
M4851 net1469 net1467 net1468 VSS nmos w=1u l=1u
M4852 net1470 net1468 VSS VSS nmos w=1u l=1u
M4853 net1469 net1467 net1471 VDD pmos w=2u l=1u
M4854 net1467 n3064 VDD VDD pmos w=2u l=1u
M4855 net1468 n3064 net1469 VDD pmos w=2u l=1u
M4856 net1468 n3065 VDD VDD pmos w=2u l=1u
M4857 n3202 net1469 VDD VDD pmos w=2u l=1u
M4858 net1471 net1468 VDD VDD pmos w=2u l=1u
M4859 n3065 n3208 VDD VDD pmos w=2u l=1u
M4860 n3065 n3208 VSS VSS nmos w=1u l=1u
M4861 n3201 n3210 net1472 VSS nmos w=1u l=1u
M4862 net1472 n3209 VSS VSS nmos w=1u l=1u
M4863 n3201 n3210 VDD VDD pmos w=2u l=1u
M4864 n3201 n3209 VDD VDD pmos w=2u l=1u
M4865 net1473 n3208 VSS VSS nmos w=1u l=1u
M4866 net1474 n3064 VSS VSS nmos w=1u l=1u
M4867 n3210 net1475 VSS VSS nmos w=1u l=1u
M4868 net1475 n3208 net1476 VSS nmos w=1u l=1u
M4869 net1475 net1473 net1474 VSS nmos w=1u l=1u
M4870 net1476 net1474 VSS VSS nmos w=1u l=1u
M4871 net1475 net1473 net1477 VDD pmos w=2u l=1u
M4872 net1473 n3208 VDD VDD pmos w=2u l=1u
M4873 net1474 n3208 net1475 VDD pmos w=2u l=1u
M4874 net1474 n3064 VDD VDD pmos w=2u l=1u
M4875 n3210 net1475 VDD VDD pmos w=2u l=1u
M4876 net1477 net1474 VDD VDD pmos w=2u l=1u
M4877 n3208 N409 net1478 VSS nmos w=1u l=1u
M4878 net1478 N171 VSS VSS nmos w=1u l=1u
M4879 n3208 N409 VDD VDD pmos w=2u l=1u
M4880 n3208 N171 VDD VDD pmos w=2u l=1u
M4881 n3064 n3063 net1479 VSS nmos w=1u l=1u
M4882 net1479 n3211 VSS VSS nmos w=1u l=1u
M4883 n3064 n3063 VDD VDD pmos w=2u l=1u
M4884 n3064 n3211 VDD VDD pmos w=2u l=1u
M4885 n3063 n3213 net1480 VSS nmos w=1u l=1u
M4886 net1480 n3212 VSS VSS nmos w=1u l=1u
M4887 n3063 n3213 VDD VDD pmos w=2u l=1u
M4888 n3063 n3212 VDD VDD pmos w=2u l=1u
M4889 n3213 n3215 net1481 VSS nmos w=1u l=1u
M4890 net1481 n3214 VSS VSS nmos w=1u l=1u
M4891 n3213 n3215 VDD VDD pmos w=2u l=1u
M4892 n3213 n3214 VDD VDD pmos w=2u l=1u
M4893 n3214 net1482 VSS VSS nmos w=1u l=1u
M4894 net1482 n3216 VSS VSS nmos w=1u l=1u
M4895 net1482 n3217 VSS VSS nmos w=1u l=1u
M4896 net1482 n3217 net1483 VDD pmos w=2u l=1u
M4897 n3214 net1482 VDD VDD pmos w=2u l=1u
M4898 net1483 n3216 VDD VDD pmos w=2u l=1u
M4899 net1484 n3074 VSS VSS nmos w=1u l=1u
M4900 net1485 n3075 VSS VSS nmos w=1u l=1u
M4901 n3212 net1486 VSS VSS nmos w=1u l=1u
M4902 net1486 n3074 net1487 VSS nmos w=1u l=1u
M4903 net1486 net1484 net1485 VSS nmos w=1u l=1u
M4904 net1487 net1485 VSS VSS nmos w=1u l=1u
M4905 net1486 net1484 net1488 VDD pmos w=2u l=1u
M4906 net1484 n3074 VDD VDD pmos w=2u l=1u
M4907 net1485 n3074 net1486 VDD pmos w=2u l=1u
M4908 net1485 n3075 VDD VDD pmos w=2u l=1u
M4909 n3212 net1486 VDD VDD pmos w=2u l=1u
M4910 net1488 net1485 VDD VDD pmos w=2u l=1u
M4911 n3075 n3218 VDD VDD pmos w=2u l=1u
M4912 n3075 n3218 VSS VSS nmos w=1u l=1u
M4913 n3211 n3220 net1489 VSS nmos w=1u l=1u
M4914 net1489 n3219 VSS VSS nmos w=1u l=1u
M4915 n3211 n3220 VDD VDD pmos w=2u l=1u
M4916 n3211 n3219 VDD VDD pmos w=2u l=1u
M4917 net1490 n3218 VSS VSS nmos w=1u l=1u
M4918 net1491 n3074 VSS VSS nmos w=1u l=1u
M4919 n3220 net1492 VSS VSS nmos w=1u l=1u
M4920 net1492 n3218 net1493 VSS nmos w=1u l=1u
M4921 net1492 net1490 net1491 VSS nmos w=1u l=1u
M4922 net1493 net1491 VSS VSS nmos w=1u l=1u
M4923 net1492 net1490 net1494 VDD pmos w=2u l=1u
M4924 net1490 n3218 VDD VDD pmos w=2u l=1u
M4925 net1491 n3218 net1492 VDD pmos w=2u l=1u
M4926 net1491 n3074 VDD VDD pmos w=2u l=1u
M4927 n3220 net1492 VDD VDD pmos w=2u l=1u
M4928 net1494 net1491 VDD VDD pmos w=2u l=1u
M4929 n3218 N392 net1495 VSS nmos w=1u l=1u
M4930 net1495 N188 VSS VSS nmos w=1u l=1u
M4931 n3218 N392 VDD VDD pmos w=2u l=1u
M4932 n3218 N188 VDD VDD pmos w=2u l=1u
M4933 n3074 n3073 net1496 VSS nmos w=1u l=1u
M4934 net1496 n3221 VSS VSS nmos w=1u l=1u
M4935 n3074 n3073 VDD VDD pmos w=2u l=1u
M4936 n3074 n3221 VDD VDD pmos w=2u l=1u
M4937 n3073 n3223 net1497 VSS nmos w=1u l=1u
M4938 net1497 n3222 VSS VSS nmos w=1u l=1u
M4939 n3073 n3223 VDD VDD pmos w=2u l=1u
M4940 n3073 n3222 VDD VDD pmos w=2u l=1u
M4941 n3223 n3225 net1498 VSS nmos w=1u l=1u
M4942 net1498 n3224 VSS VSS nmos w=1u l=1u
M4943 n3223 n3225 VDD VDD pmos w=2u l=1u
M4944 n3223 n3224 VDD VDD pmos w=2u l=1u
M4945 n3224 net1499 VSS VSS nmos w=1u l=1u
M4946 net1499 n3226 VSS VSS nmos w=1u l=1u
M4947 net1499 n3227 VSS VSS nmos w=1u l=1u
M4948 net1499 n3227 net1500 VDD pmos w=2u l=1u
M4949 n3224 net1499 VDD VDD pmos w=2u l=1u
M4950 net1500 n3226 VDD VDD pmos w=2u l=1u
M4951 net1501 n3084 VSS VSS nmos w=1u l=1u
M4952 net1502 n3085 VSS VSS nmos w=1u l=1u
M4953 n3222 net1503 VSS VSS nmos w=1u l=1u
M4954 net1503 n3084 net1504 VSS nmos w=1u l=1u
M4955 net1503 net1501 net1502 VSS nmos w=1u l=1u
M4956 net1504 net1502 VSS VSS nmos w=1u l=1u
M4957 net1503 net1501 net1505 VDD pmos w=2u l=1u
M4958 net1501 n3084 VDD VDD pmos w=2u l=1u
M4959 net1502 n3084 net1503 VDD pmos w=2u l=1u
M4960 net1502 n3085 VDD VDD pmos w=2u l=1u
M4961 n3222 net1503 VDD VDD pmos w=2u l=1u
M4962 net1505 net1502 VDD VDD pmos w=2u l=1u
M4963 n3085 n3228 VDD VDD pmos w=2u l=1u
M4964 n3085 n3228 VSS VSS nmos w=1u l=1u
M4965 n3221 n3230 net1506 VSS nmos w=1u l=1u
M4966 net1506 n3229 VSS VSS nmos w=1u l=1u
M4967 n3221 n3230 VDD VDD pmos w=2u l=1u
M4968 n3221 n3229 VDD VDD pmos w=2u l=1u
M4969 net1507 n3228 VSS VSS nmos w=1u l=1u
M4970 net1508 n3084 VSS VSS nmos w=1u l=1u
M4971 n3230 net1509 VSS VSS nmos w=1u l=1u
M4972 net1509 n3228 net1510 VSS nmos w=1u l=1u
M4973 net1509 net1507 net1508 VSS nmos w=1u l=1u
M4974 net1510 net1508 VSS VSS nmos w=1u l=1u
M4975 net1509 net1507 net1511 VDD pmos w=2u l=1u
M4976 net1507 n3228 VDD VDD pmos w=2u l=1u
M4977 net1508 n3228 net1509 VDD pmos w=2u l=1u
M4978 net1508 n3084 VDD VDD pmos w=2u l=1u
M4979 n3230 net1509 VDD VDD pmos w=2u l=1u
M4980 net1511 net1508 VDD VDD pmos w=2u l=1u
M4981 n3228 N375 net1512 VSS nmos w=1u l=1u
M4982 net1512 N205 VSS VSS nmos w=1u l=1u
M4983 n3228 N375 VDD VDD pmos w=2u l=1u
M4984 n3228 N205 VDD VDD pmos w=2u l=1u
M4985 n3084 n3083 net1513 VSS nmos w=1u l=1u
M4986 net1513 n3231 VSS VSS nmos w=1u l=1u
M4987 n3084 n3083 VDD VDD pmos w=2u l=1u
M4988 n3084 n3231 VDD VDD pmos w=2u l=1u
M4989 n3083 n3233 net1514 VSS nmos w=1u l=1u
M4990 net1514 n3232 VSS VSS nmos w=1u l=1u
M4991 n3083 n3233 VDD VDD pmos w=2u l=1u
M4992 n3083 n3232 VDD VDD pmos w=2u l=1u
M4993 n3233 n3235 net1515 VSS nmos w=1u l=1u
M4994 net1515 n3234 VSS VSS nmos w=1u l=1u
M4995 n3233 n3235 VDD VDD pmos w=2u l=1u
M4996 n3233 n3234 VDD VDD pmos w=2u l=1u
M4997 n3234 net1516 VSS VSS nmos w=1u l=1u
M4998 net1516 n3236 VSS VSS nmos w=1u l=1u
M4999 net1516 n3237 VSS VSS nmos w=1u l=1u
M5000 net1516 n3237 net1517 VDD pmos w=2u l=1u
M5001 n3234 net1516 VDD VDD pmos w=2u l=1u
M5002 net1517 n3236 VDD VDD pmos w=2u l=1u
M5003 net1518 n3095 VSS VSS nmos w=1u l=1u
M5004 net1519 n3096 VSS VSS nmos w=1u l=1u
M5005 n3232 net1520 VSS VSS nmos w=1u l=1u
M5006 net1520 n3095 net1521 VSS nmos w=1u l=1u
M5007 net1520 net1518 net1519 VSS nmos w=1u l=1u
M5008 net1521 net1519 VSS VSS nmos w=1u l=1u
M5009 net1520 net1518 net1522 VDD pmos w=2u l=1u
M5010 net1518 n3095 VDD VDD pmos w=2u l=1u
M5011 net1519 n3095 net1520 VDD pmos w=2u l=1u
M5012 net1519 n3096 VDD VDD pmos w=2u l=1u
M5013 n3232 net1520 VDD VDD pmos w=2u l=1u
M5014 net1522 net1519 VDD VDD pmos w=2u l=1u
M5015 n3095 n3238 VDD VDD pmos w=2u l=1u
M5016 n3095 n3238 VSS VSS nmos w=1u l=1u
M5017 n3231 n3240 net1523 VSS nmos w=1u l=1u
M5018 net1523 n3239 VSS VSS nmos w=1u l=1u
M5019 n3231 n3240 VDD VDD pmos w=2u l=1u
M5020 n3231 n3239 VDD VDD pmos w=2u l=1u
M5021 net1524 n3096 VSS VSS nmos w=1u l=1u
M5022 net1525 n3238 VSS VSS nmos w=1u l=1u
M5023 n3240 net1526 VSS VSS nmos w=1u l=1u
M5024 net1526 n3096 net1527 VSS nmos w=1u l=1u
M5025 net1526 net1524 net1525 VSS nmos w=1u l=1u
M5026 net1527 net1525 VSS VSS nmos w=1u l=1u
M5027 net1526 net1524 net1528 VDD pmos w=2u l=1u
M5028 net1524 n3096 VDD VDD pmos w=2u l=1u
M5029 net1525 n3096 net1526 VDD pmos w=2u l=1u
M5030 net1525 n3238 VDD VDD pmos w=2u l=1u
M5031 n3240 net1526 VDD VDD pmos w=2u l=1u
M5032 net1528 net1525 VDD VDD pmos w=2u l=1u
M5033 n3096 N358 net1529 VSS nmos w=1u l=1u
M5034 net1529 N222 VSS VSS nmos w=1u l=1u
M5035 n3096 N358 VDD VDD pmos w=2u l=1u
M5036 n3096 N222 VDD VDD pmos w=2u l=1u
M5037 n3238 n3093 net1530 VSS nmos w=1u l=1u
M5038 net1530 n3241 VSS VSS nmos w=1u l=1u
M5039 n3238 n3093 VDD VDD pmos w=2u l=1u
M5040 n3238 n3241 VDD VDD pmos w=2u l=1u
M5041 n3093 n3243 net1531 VSS nmos w=1u l=1u
M5042 net1531 n3242 VSS VSS nmos w=1u l=1u
M5043 n3093 n3243 VDD VDD pmos w=2u l=1u
M5044 n3093 n3242 VDD VDD pmos w=2u l=1u
M5045 n3243 n3245 net1532 VSS nmos w=1u l=1u
M5046 net1532 n3244 VSS VSS nmos w=1u l=1u
M5047 n3243 n3245 VDD VDD pmos w=2u l=1u
M5048 n3243 n3244 VDD VDD pmos w=2u l=1u
M5049 n3241 n3244 net1533 VSS nmos w=1u l=1u
M5050 net1533 n3246 VSS VSS nmos w=1u l=1u
M5051 n3241 n3244 VDD VDD pmos w=2u l=1u
M5052 n3241 n3246 VDD VDD pmos w=2u l=1u
M5053 n3244 n3248 net1534 VSS nmos w=1u l=1u
M5054 net1534 n3247 VSS VSS nmos w=1u l=1u
M5055 n3244 n3248 VDD VDD pmos w=2u l=1u
M5056 n3244 n3247 VDD VDD pmos w=2u l=1u
M5057 n3246 n3242 VSS VSS nmos w=1u l=1u
M5058 n3246 n3249 VSS VSS nmos w=1u l=1u
M5059 n3246 n3242 net1535 VDD pmos w=2u l=1u
M5060 net1535 n3249 VDD VDD pmos w=2u l=1u
M5061 n3242 net1536 VSS VSS nmos w=1u l=1u
M5062 net1537 n3250 VSS VSS nmos w=1u l=1u
M5063 net1536 n3108 net1537 VSS nmos w=1u l=1u
M5064 net1536 n3250 VDD VDD pmos w=2u l=1u
M5065 net1536 n3108 VDD VDD pmos w=2u l=1u
M5066 n3242 net1536 VDD VDD pmos w=2u l=1u
M5067 n3250 N341 net1538 VSS nmos w=1u l=1u
M5068 net1538 n3251 VSS VSS nmos w=1u l=1u
M5069 n3250 N341 VDD VDD pmos w=2u l=1u
M5070 n3250 n3251 VDD VDD pmos w=2u l=1u
M5071 n3251 n3253 VSS VSS nmos w=1u l=1u
M5072 n3251 n3252 VSS VSS nmos w=1u l=1u
M5073 n3251 n3253 net1539 VDD pmos w=2u l=1u
M5074 net1539 n3252 VDD VDD pmos w=2u l=1u
M5075 n3253 n3255 VSS VSS nmos w=1u l=1u
M5076 n3253 n3254 VSS VSS nmos w=1u l=1u
M5077 n3253 n3255 net1540 VDD pmos w=2u l=1u
M5078 net1540 n3254 VDD VDD pmos w=2u l=1u
M5079 n3255 n2270 net1541 VSS nmos w=1u l=1u
M5080 net1541 n3256 VSS VSS nmos w=1u l=1u
M5081 n3255 n2270 VDD VDD pmos w=2u l=1u
M5082 n3255 n3256 VDD VDD pmos w=2u l=1u
M5083 n3256 n3257 net1542 VSS nmos w=1u l=1u
M5084 net1542 N239 VSS VSS nmos w=1u l=1u
M5085 n3256 n3257 VDD VDD pmos w=2u l=1u
M5086 n3256 N239 VDD VDD pmos w=2u l=1u
M5087 n3254 n3111 VDD VDD pmos w=2u l=1u
M5088 n3254 n3111 VSS VSS nmos w=1u l=1u
M5089 n3252 n3111 VSS VSS nmos w=1u l=1u
M5090 n3252 N324 VSS VSS nmos w=1u l=1u
M5091 n3252 n3111 net1543 VDD pmos w=2u l=1u
M5092 net1543 N324 VDD VDD pmos w=2u l=1u
M5093 n3108 n3259 net1544 VSS nmos w=1u l=1u
M5094 net1544 n3258 VSS VSS nmos w=1u l=1u
M5095 n3108 n3259 VDD VDD pmos w=2u l=1u
M5096 n3108 n3258 VDD VDD pmos w=2u l=1u
M5097 n3259 N239 net1545 VSS nmos w=1u l=1u
M5098 net1545 N341 VSS VSS nmos w=1u l=1u
M5099 n3259 N239 VDD VDD pmos w=2u l=1u
M5100 n3259 N341 VDD VDD pmos w=2u l=1u
M5101 net1546 n3110 VSS VSS nmos w=1u l=1u
M5102 net1547 n3111 VSS VSS nmos w=1u l=1u
M5103 n3258 net1548 VSS VSS nmos w=1u l=1u
M5104 net1548 n3110 net1549 VSS nmos w=1u l=1u
M5105 net1548 net1546 net1547 VSS nmos w=1u l=1u
M5106 net1549 net1547 VSS VSS nmos w=1u l=1u
M5107 net1548 net1546 net1550 VDD pmos w=2u l=1u
M5108 net1546 n3110 VDD VDD pmos w=2u l=1u
M5109 net1547 n3110 net1548 VDD pmos w=2u l=1u
M5110 net1547 n3111 VDD VDD pmos w=2u l=1u
M5111 n3258 net1548 VDD VDD pmos w=2u l=1u
M5112 net1550 net1547 VDD VDD pmos w=2u l=1u
M5113 n3110 N256 net1551 VSS nmos w=1u l=1u
M5114 net1551 N324 VSS VSS nmos w=1u l=1u
M5115 n3110 N256 VDD VDD pmos w=2u l=1u
M5116 n3110 N324 VDD VDD pmos w=2u l=1u
M5117 n3111 n3261 net1552 VSS nmos w=1u l=1u
M5118 net1552 n3260 VSS VSS nmos w=1u l=1u
M5119 n3111 n3261 VDD VDD pmos w=2u l=1u
M5120 n3111 n3260 VDD VDD pmos w=2u l=1u
M5121 n3261 n3263 net1553 VSS nmos w=1u l=1u
M5122 net1553 n3262 VSS VSS nmos w=1u l=1u
M5123 n3261 n3263 VDD VDD pmos w=2u l=1u
M5124 n3261 n3262 VDD VDD pmos w=2u l=1u
M5125 n3239 n3265 VSS VSS nmos w=1u l=1u
M5126 n3239 n3264 VSS VSS nmos w=1u l=1u
M5127 n3239 n3265 net1554 VDD pmos w=2u l=1u
M5128 net1554 n3264 VDD VDD pmos w=2u l=1u
M5129 n3265 n3236 VSS VSS nmos w=1u l=1u
M5130 n3265 n3237 VSS VSS nmos w=1u l=1u
M5131 n3265 n3236 net1555 VDD pmos w=2u l=1u
M5132 net1555 n3237 VDD VDD pmos w=2u l=1u
M5133 n3264 n3235 VDD VDD pmos w=2u l=1u
M5134 n3264 n3235 VSS VSS nmos w=1u l=1u
M5135 n3229 n3267 VSS VSS nmos w=1u l=1u
M5136 n3229 n3266 VSS VSS nmos w=1u l=1u
M5137 n3229 n3267 net1556 VDD pmos w=2u l=1u
M5138 net1556 n3266 VDD VDD pmos w=2u l=1u
M5139 n3267 n3226 VSS VSS nmos w=1u l=1u
M5140 n3267 n3227 VSS VSS nmos w=1u l=1u
M5141 n3267 n3226 net1557 VDD pmos w=2u l=1u
M5142 net1557 n3227 VDD VDD pmos w=2u l=1u
M5143 n3266 n3225 VDD VDD pmos w=2u l=1u
M5144 n3266 n3225 VSS VSS nmos w=1u l=1u
M5145 n3219 n3269 VSS VSS nmos w=1u l=1u
M5146 n3219 n3268 VSS VSS nmos w=1u l=1u
M5147 n3219 n3269 net1558 VDD pmos w=2u l=1u
M5148 net1558 n3268 VDD VDD pmos w=2u l=1u
M5149 n3269 n3216 VSS VSS nmos w=1u l=1u
M5150 n3269 n3217 VSS VSS nmos w=1u l=1u
M5151 n3269 n3216 net1559 VDD pmos w=2u l=1u
M5152 net1559 n3217 VDD VDD pmos w=2u l=1u
M5153 n3268 n3215 VDD VDD pmos w=2u l=1u
M5154 n3268 n3215 VSS VSS nmos w=1u l=1u
M5155 n3209 n3271 VSS VSS nmos w=1u l=1u
M5156 n3209 n3270 VSS VSS nmos w=1u l=1u
M5157 n3209 n3271 net1560 VDD pmos w=2u l=1u
M5158 net1560 n3270 VDD VDD pmos w=2u l=1u
M5159 n3271 n3206 VSS VSS nmos w=1u l=1u
M5160 n3271 n3207 VSS VSS nmos w=1u l=1u
M5161 n3271 n3206 net1561 VDD pmos w=2u l=1u
M5162 net1561 n3207 VDD VDD pmos w=2u l=1u
M5163 n3270 n3205 VDD VDD pmos w=2u l=1u
M5164 n3270 n3205 VSS VSS nmos w=1u l=1u
M5165 n3199 n3273 VSS VSS nmos w=1u l=1u
M5166 n3199 n3272 VSS VSS nmos w=1u l=1u
M5167 n3199 n3273 net1562 VDD pmos w=2u l=1u
M5168 net1562 n3272 VDD VDD pmos w=2u l=1u
M5169 n3273 n3196 VSS VSS nmos w=1u l=1u
M5170 n3273 n3197 VSS VSS nmos w=1u l=1u
M5171 n3273 n3196 net1563 VDD pmos w=2u l=1u
M5172 net1563 n3197 VDD VDD pmos w=2u l=1u
M5173 n3272 n3195 VDD VDD pmos w=2u l=1u
M5174 n3272 n3195 VSS VSS nmos w=1u l=1u
M5175 n3189 n3275 VSS VSS nmos w=1u l=1u
M5176 n3189 n3274 VSS VSS nmos w=1u l=1u
M5177 n3189 n3275 net1564 VDD pmos w=2u l=1u
M5178 net1564 n3274 VDD VDD pmos w=2u l=1u
M5179 n3275 n3186 VSS VSS nmos w=1u l=1u
M5180 n3275 n3187 VSS VSS nmos w=1u l=1u
M5181 n3275 n3186 net1565 VDD pmos w=2u l=1u
M5182 net1565 n3187 VDD VDD pmos w=2u l=1u
M5183 n3274 n3185 VDD VDD pmos w=2u l=1u
M5184 n3274 n3185 VSS VSS nmos w=1u l=1u
M5185 n3179 n3277 VSS VSS nmos w=1u l=1u
M5186 n3179 n3276 VSS VSS nmos w=1u l=1u
M5187 n3179 n3277 net1566 VDD pmos w=2u l=1u
M5188 net1566 n3276 VDD VDD pmos w=2u l=1u
M5189 n3277 n3176 VSS VSS nmos w=1u l=1u
M5190 n3277 n3177 VSS VSS nmos w=1u l=1u
M5191 n3277 n3176 net1567 VDD pmos w=2u l=1u
M5192 net1567 n3177 VDD VDD pmos w=2u l=1u
M5193 n3276 n3175 VDD VDD pmos w=2u l=1u
M5194 n3276 n3175 VSS VSS nmos w=1u l=1u
M5195 n3169 n3279 VSS VSS nmos w=1u l=1u
M5196 n3169 n3278 VSS VSS nmos w=1u l=1u
M5197 n3169 n3279 net1568 VDD pmos w=2u l=1u
M5198 net1568 n3278 VDD VDD pmos w=2u l=1u
M5199 n3279 n3166 VSS VSS nmos w=1u l=1u
M5200 n3279 n3167 VSS VSS nmos w=1u l=1u
M5201 n3279 n3166 net1569 VDD pmos w=2u l=1u
M5202 net1569 n3167 VDD VDD pmos w=2u l=1u
M5203 n3278 n3165 VDD VDD pmos w=2u l=1u
M5204 n3278 n3165 VSS VSS nmos w=1u l=1u
M5205 n3159 n3281 VSS VSS nmos w=1u l=1u
M5206 n3159 n3280 VSS VSS nmos w=1u l=1u
M5207 n3159 n3281 net1570 VDD pmos w=2u l=1u
M5208 net1570 n3280 VDD VDD pmos w=2u l=1u
M5209 n3281 n3156 VSS VSS nmos w=1u l=1u
M5210 n3281 n3157 VSS VSS nmos w=1u l=1u
M5211 n3281 n3156 net1571 VDD pmos w=2u l=1u
M5212 net1571 n3157 VDD VDD pmos w=2u l=1u
M5213 n3280 n3155 VDD VDD pmos w=2u l=1u
M5214 n3280 n3155 VSS VSS nmos w=1u l=1u
M5215 n3149 n3283 VSS VSS nmos w=1u l=1u
M5216 n3149 n3282 VSS VSS nmos w=1u l=1u
M5217 n3149 n3283 net1572 VDD pmos w=2u l=1u
M5218 net1572 n3282 VDD VDD pmos w=2u l=1u
M5219 n3283 n3146 VSS VSS nmos w=1u l=1u
M5220 n3283 n3147 VSS VSS nmos w=1u l=1u
M5221 n3283 n3146 net1573 VDD pmos w=2u l=1u
M5222 net1573 n3147 VDD VDD pmos w=2u l=1u
M5223 n3282 n3145 VDD VDD pmos w=2u l=1u
M5224 n3282 n3145 VSS VSS nmos w=1u l=1u
M5225 n2998 N528 net1574 VSS nmos w=1u l=1u
M5226 net1574 N52 VSS VSS nmos w=1u l=1u
M5227 n2998 N528 VDD VDD pmos w=2u l=1u
M5228 n2998 N52 VDD VDD pmos w=2u l=1u
M5229 N6160 n3284 net1575 VSS nmos w=1u l=1u
M5230 net1575 n3134 VSS VSS nmos w=1u l=1u
M5231 N6160 n3284 VDD VDD pmos w=2u l=1u
M5232 N6160 n3134 VDD VDD pmos w=2u l=1u
M5233 n3284 net1576 VSS VSS nmos w=1u l=1u
M5234 net1576 n3285 VSS VSS nmos w=1u l=1u
M5235 net1576 n3286 VSS VSS nmos w=1u l=1u
M5236 net1576 n3286 net1577 VDD pmos w=2u l=1u
M5237 n3284 net1576 VDD VDD pmos w=2u l=1u
M5238 net1577 n3285 VDD VDD pmos w=2u l=1u
M5239 n3134 n3286 net1578 VSS nmos w=1u l=1u
M5240 net1578 n3285 VSS VSS nmos w=1u l=1u
M5241 n3134 n3286 VDD VDD pmos w=2u l=1u
M5242 n3134 n3285 VDD VDD pmos w=2u l=1u
M5243 net1579 n3136 VSS VSS nmos w=1u l=1u
M5244 net1580 n3135 VSS VSS nmos w=1u l=1u
M5245 n3285 net1581 VSS VSS nmos w=1u l=1u
M5246 net1581 n3136 net1582 VSS nmos w=1u l=1u
M5247 net1581 net1579 net1580 VSS nmos w=1u l=1u
M5248 net1582 net1580 VSS VSS nmos w=1u l=1u
M5249 net1581 net1579 net1583 VDD pmos w=2u l=1u
M5250 net1579 n3136 VDD VDD pmos w=2u l=1u
M5251 net1580 n3136 net1581 VDD pmos w=2u l=1u
M5252 net1580 n3135 VDD VDD pmos w=2u l=1u
M5253 n3285 net1581 VDD VDD pmos w=2u l=1u
M5254 net1583 net1580 VDD VDD pmos w=2u l=1u
M5255 n3136 n3288 net1584 VSS nmos w=1u l=1u
M5256 net1584 n3287 VSS VSS nmos w=1u l=1u
M5257 n3136 n3288 VDD VDD pmos w=2u l=1u
M5258 n3136 n3287 VDD VDD pmos w=2u l=1u
M5259 n3287 n3290 net1585 VSS nmos w=1u l=1u
M5260 net1585 n3289 VSS VSS nmos w=1u l=1u
M5261 n3287 n3290 VDD VDD pmos w=2u l=1u
M5262 n3287 n3289 VDD VDD pmos w=2u l=1u
M5263 n3290 N528 net1586 VSS nmos w=1u l=1u
M5264 net1586 N18 VSS VSS nmos w=1u l=1u
M5265 n3290 N528 VDD VDD pmos w=2u l=1u
M5266 n3290 N18 VDD VDD pmos w=2u l=1u
M5267 net1587 n3139 VSS VSS nmos w=1u l=1u
M5268 net1588 n3140 VSS VSS nmos w=1u l=1u
M5269 n3135 net1589 VSS VSS nmos w=1u l=1u
M5270 net1589 n3139 net1590 VSS nmos w=1u l=1u
M5271 net1589 net1587 net1588 VSS nmos w=1u l=1u
M5272 net1590 net1588 VSS VSS nmos w=1u l=1u
M5273 net1589 net1587 net1591 VDD pmos w=2u l=1u
M5274 net1587 n3139 VDD VDD pmos w=2u l=1u
M5275 net1588 n3139 net1589 VDD pmos w=2u l=1u
M5276 net1588 n3140 VDD VDD pmos w=2u l=1u
M5277 n3135 net1589 VDD VDD pmos w=2u l=1u
M5278 net1591 net1588 VDD VDD pmos w=2u l=1u
M5279 n3139 net1592 VSS VSS nmos w=1u l=1u
M5280 net1593 n3138 VSS VSS nmos w=1u l=1u
M5281 net1592 n3291 net1593 VSS nmos w=1u l=1u
M5282 net1592 n3138 VDD VDD pmos w=2u l=1u
M5283 net1592 n3291 VDD VDD pmos w=2u l=1u
M5284 n3139 net1592 VDD VDD pmos w=2u l=1u
M5285 n3138 n3293 net1594 VSS nmos w=1u l=1u
M5286 net1594 n3292 VSS VSS nmos w=1u l=1u
M5287 n3138 n3293 VDD VDD pmos w=2u l=1u
M5288 n3138 n3292 VDD VDD pmos w=2u l=1u
M5289 n3293 n3295 net1595 VSS nmos w=1u l=1u
M5290 net1595 n3294 VSS VSS nmos w=1u l=1u
M5291 n3293 n3295 VDD VDD pmos w=2u l=1u
M5292 n3293 n3294 VDD VDD pmos w=2u l=1u
M5293 n3294 net1596 VSS VSS nmos w=1u l=1u
M5294 net1596 n3296 VSS VSS nmos w=1u l=1u
M5295 net1596 n3297 VSS VSS nmos w=1u l=1u
M5296 net1596 n3297 net1597 VDD pmos w=2u l=1u
M5297 n3294 net1596 VDD VDD pmos w=2u l=1u
M5298 net1597 n3296 VDD VDD pmos w=2u l=1u
M5299 net1598 n3146 VSS VSS nmos w=1u l=1u
M5300 net1599 n3147 VSS VSS nmos w=1u l=1u
M5301 n3292 net1600 VSS VSS nmos w=1u l=1u
M5302 net1600 n3146 net1601 VSS nmos w=1u l=1u
M5303 net1600 net1598 net1599 VSS nmos w=1u l=1u
M5304 net1601 net1599 VSS VSS nmos w=1u l=1u
M5305 net1600 net1598 net1602 VDD pmos w=2u l=1u
M5306 net1598 n3146 VDD VDD pmos w=2u l=1u
M5307 net1599 n3146 net1600 VDD pmos w=2u l=1u
M5308 net1599 n3147 VDD VDD pmos w=2u l=1u
M5309 n3292 net1600 VDD VDD pmos w=2u l=1u
M5310 net1602 net1599 VDD VDD pmos w=2u l=1u
M5311 n3147 n3298 VDD VDD pmos w=2u l=1u
M5312 n3147 n3298 VSS VSS nmos w=1u l=1u
M5313 n3291 n3300 net1603 VSS nmos w=1u l=1u
M5314 net1603 n3299 VSS VSS nmos w=1u l=1u
M5315 n3291 n3300 VDD VDD pmos w=2u l=1u
M5316 n3291 n3299 VDD VDD pmos w=2u l=1u
M5317 net1604 n3298 VSS VSS nmos w=1u l=1u
M5318 net1605 n3146 VSS VSS nmos w=1u l=1u
M5319 n3300 net1606 VSS VSS nmos w=1u l=1u
M5320 net1606 n3298 net1607 VSS nmos w=1u l=1u
M5321 net1606 net1604 net1605 VSS nmos w=1u l=1u
M5322 net1607 net1605 VSS VSS nmos w=1u l=1u
M5323 net1606 net1604 net1608 VDD pmos w=2u l=1u
M5324 net1604 n3298 VDD VDD pmos w=2u l=1u
M5325 net1605 n3298 net1606 VDD pmos w=2u l=1u
M5326 net1605 n3146 VDD VDD pmos w=2u l=1u
M5327 n3300 net1606 VDD VDD pmos w=2u l=1u
M5328 net1608 net1605 VDD VDD pmos w=2u l=1u
M5329 n3298 N511 net1609 VSS nmos w=1u l=1u
M5330 net1609 N52 VSS VSS nmos w=1u l=1u
M5331 n3298 N511 VDD VDD pmos w=2u l=1u
M5332 n3298 N52 VDD VDD pmos w=2u l=1u
M5333 n3146 n3145 net1610 VSS nmos w=1u l=1u
M5334 net1610 n3301 VSS VSS nmos w=1u l=1u
M5335 n3146 n3145 VDD VDD pmos w=2u l=1u
M5336 n3146 n3301 VDD VDD pmos w=2u l=1u
M5337 n3145 n3303 net1611 VSS nmos w=1u l=1u
M5338 net1611 n3302 VSS VSS nmos w=1u l=1u
M5339 n3145 n3303 VDD VDD pmos w=2u l=1u
M5340 n3145 n3302 VDD VDD pmos w=2u l=1u
M5341 n3303 n3305 net1612 VSS nmos w=1u l=1u
M5342 net1612 n3304 VSS VSS nmos w=1u l=1u
M5343 n3303 n3305 VDD VDD pmos w=2u l=1u
M5344 n3303 n3304 VDD VDD pmos w=2u l=1u
M5345 n3304 net1613 VSS VSS nmos w=1u l=1u
M5346 net1613 n3306 VSS VSS nmos w=1u l=1u
M5347 net1613 n3307 VSS VSS nmos w=1u l=1u
M5348 net1613 n3307 net1614 VDD pmos w=2u l=1u
M5349 n3304 net1613 VDD VDD pmos w=2u l=1u
M5350 net1614 n3306 VDD VDD pmos w=2u l=1u
M5351 net1615 n3156 VSS VSS nmos w=1u l=1u
M5352 net1616 n3157 VSS VSS nmos w=1u l=1u
M5353 n3302 net1617 VSS VSS nmos w=1u l=1u
M5354 net1617 n3156 net1618 VSS nmos w=1u l=1u
M5355 net1617 net1615 net1616 VSS nmos w=1u l=1u
M5356 net1618 net1616 VSS VSS nmos w=1u l=1u
M5357 net1617 net1615 net1619 VDD pmos w=2u l=1u
M5358 net1615 n3156 VDD VDD pmos w=2u l=1u
M5359 net1616 n3156 net1617 VDD pmos w=2u l=1u
M5360 net1616 n3157 VDD VDD pmos w=2u l=1u
M5361 n3302 net1617 VDD VDD pmos w=2u l=1u
M5362 net1619 net1616 VDD VDD pmos w=2u l=1u
M5363 n3157 n3308 VDD VDD pmos w=2u l=1u
M5364 n3157 n3308 VSS VSS nmos w=1u l=1u
M5365 n3301 n3310 net1620 VSS nmos w=1u l=1u
M5366 net1620 n3309 VSS VSS nmos w=1u l=1u
M5367 n3301 n3310 VDD VDD pmos w=2u l=1u
M5368 n3301 n3309 VDD VDD pmos w=2u l=1u
M5369 net1621 n3308 VSS VSS nmos w=1u l=1u
M5370 net1622 n3156 VSS VSS nmos w=1u l=1u
M5371 n3310 net1623 VSS VSS nmos w=1u l=1u
M5372 net1623 n3308 net1624 VSS nmos w=1u l=1u
M5373 net1623 net1621 net1622 VSS nmos w=1u l=1u
M5374 net1624 net1622 VSS VSS nmos w=1u l=1u
M5375 net1623 net1621 net1625 VDD pmos w=2u l=1u
M5376 net1621 n3308 VDD VDD pmos w=2u l=1u
M5377 net1622 n3308 net1623 VDD pmos w=2u l=1u
M5378 net1622 n3156 VDD VDD pmos w=2u l=1u
M5379 n3310 net1623 VDD VDD pmos w=2u l=1u
M5380 net1625 net1622 VDD VDD pmos w=2u l=1u
M5381 n3308 N494 net1626 VSS nmos w=1u l=1u
M5382 net1626 N69 VSS VSS nmos w=1u l=1u
M5383 n3308 N494 VDD VDD pmos w=2u l=1u
M5384 n3308 N69 VDD VDD pmos w=2u l=1u
M5385 n3156 n3155 net1627 VSS nmos w=1u l=1u
M5386 net1627 n3311 VSS VSS nmos w=1u l=1u
M5387 n3156 n3155 VDD VDD pmos w=2u l=1u
M5388 n3156 n3311 VDD VDD pmos w=2u l=1u
M5389 n3155 n3313 net1628 VSS nmos w=1u l=1u
M5390 net1628 n3312 VSS VSS nmos w=1u l=1u
M5391 n3155 n3313 VDD VDD pmos w=2u l=1u
M5392 n3155 n3312 VDD VDD pmos w=2u l=1u
M5393 n3313 n3315 net1629 VSS nmos w=1u l=1u
M5394 net1629 n3314 VSS VSS nmos w=1u l=1u
M5395 n3313 n3315 VDD VDD pmos w=2u l=1u
M5396 n3313 n3314 VDD VDD pmos w=2u l=1u
M5397 n3314 net1630 VSS VSS nmos w=1u l=1u
M5398 net1630 n3316 VSS VSS nmos w=1u l=1u
M5399 net1630 n3317 VSS VSS nmos w=1u l=1u
M5400 net1630 n3317 net1631 VDD pmos w=2u l=1u
M5401 n3314 net1630 VDD VDD pmos w=2u l=1u
M5402 net1631 n3316 VDD VDD pmos w=2u l=1u
M5403 net1632 n3166 VSS VSS nmos w=1u l=1u
M5404 net1633 n3167 VSS VSS nmos w=1u l=1u
M5405 n3312 net1634 VSS VSS nmos w=1u l=1u
M5406 net1634 n3166 net1635 VSS nmos w=1u l=1u
M5407 net1634 net1632 net1633 VSS nmos w=1u l=1u
M5408 net1635 net1633 VSS VSS nmos w=1u l=1u
M5409 net1634 net1632 net1636 VDD pmos w=2u l=1u
M5410 net1632 n3166 VDD VDD pmos w=2u l=1u
M5411 net1633 n3166 net1634 VDD pmos w=2u l=1u
M5412 net1633 n3167 VDD VDD pmos w=2u l=1u
M5413 n3312 net1634 VDD VDD pmos w=2u l=1u
M5414 net1636 net1633 VDD VDD pmos w=2u l=1u
M5415 n3167 n3318 VDD VDD pmos w=2u l=1u
M5416 n3167 n3318 VSS VSS nmos w=1u l=1u
M5417 n3311 n3320 net1637 VSS nmos w=1u l=1u
M5418 net1637 n3319 VSS VSS nmos w=1u l=1u
M5419 n3311 n3320 VDD VDD pmos w=2u l=1u
M5420 n3311 n3319 VDD VDD pmos w=2u l=1u
M5421 net1638 n3318 VSS VSS nmos w=1u l=1u
M5422 net1639 n3166 VSS VSS nmos w=1u l=1u
M5423 n3320 net1640 VSS VSS nmos w=1u l=1u
M5424 net1640 n3318 net1641 VSS nmos w=1u l=1u
M5425 net1640 net1638 net1639 VSS nmos w=1u l=1u
M5426 net1641 net1639 VSS VSS nmos w=1u l=1u
M5427 net1640 net1638 net1642 VDD pmos w=2u l=1u
M5428 net1638 n3318 VDD VDD pmos w=2u l=1u
M5429 net1639 n3318 net1640 VDD pmos w=2u l=1u
M5430 net1639 n3166 VDD VDD pmos w=2u l=1u
M5431 n3320 net1640 VDD VDD pmos w=2u l=1u
M5432 net1642 net1639 VDD VDD pmos w=2u l=1u
M5433 n3318 N477 net1643 VSS nmos w=1u l=1u
M5434 net1643 N86 VSS VSS nmos w=1u l=1u
M5435 n3318 N477 VDD VDD pmos w=2u l=1u
M5436 n3318 N86 VDD VDD pmos w=2u l=1u
M5437 n3166 n3165 net1644 VSS nmos w=1u l=1u
M5438 net1644 n3321 VSS VSS nmos w=1u l=1u
M5439 n3166 n3165 VDD VDD pmos w=2u l=1u
M5440 n3166 n3321 VDD VDD pmos w=2u l=1u
M5441 n3165 n3323 net1645 VSS nmos w=1u l=1u
M5442 net1645 n3322 VSS VSS nmos w=1u l=1u
M5443 n3165 n3323 VDD VDD pmos w=2u l=1u
M5444 n3165 n3322 VDD VDD pmos w=2u l=1u
M5445 n3323 n3325 net1646 VSS nmos w=1u l=1u
M5446 net1646 n3324 VSS VSS nmos w=1u l=1u
M5447 n3323 n3325 VDD VDD pmos w=2u l=1u
M5448 n3323 n3324 VDD VDD pmos w=2u l=1u
M5449 n3324 net1647 VSS VSS nmos w=1u l=1u
M5450 net1647 n3326 VSS VSS nmos w=1u l=1u
M5451 net1647 n3327 VSS VSS nmos w=1u l=1u
M5452 net1647 n3327 net1648 VDD pmos w=2u l=1u
M5453 n3324 net1647 VDD VDD pmos w=2u l=1u
M5454 net1648 n3326 VDD VDD pmos w=2u l=1u
M5455 net1649 n3176 VSS VSS nmos w=1u l=1u
M5456 net1650 n3177 VSS VSS nmos w=1u l=1u
M5457 n3322 net1651 VSS VSS nmos w=1u l=1u
M5458 net1651 n3176 net1652 VSS nmos w=1u l=1u
M5459 net1651 net1649 net1650 VSS nmos w=1u l=1u
M5460 net1652 net1650 VSS VSS nmos w=1u l=1u
M5461 net1651 net1649 net1653 VDD pmos w=2u l=1u
M5462 net1649 n3176 VDD VDD pmos w=2u l=1u
M5463 net1650 n3176 net1651 VDD pmos w=2u l=1u
M5464 net1650 n3177 VDD VDD pmos w=2u l=1u
M5465 n3322 net1651 VDD VDD pmos w=2u l=1u
M5466 net1653 net1650 VDD VDD pmos w=2u l=1u
M5467 n3177 n3328 VDD VDD pmos w=2u l=1u
M5468 n3177 n3328 VSS VSS nmos w=1u l=1u
M5469 n3321 n3330 net1654 VSS nmos w=1u l=1u
M5470 net1654 n3329 VSS VSS nmos w=1u l=1u
M5471 n3321 n3330 VDD VDD pmos w=2u l=1u
M5472 n3321 n3329 VDD VDD pmos w=2u l=1u
M5473 net1655 n3328 VSS VSS nmos w=1u l=1u
M5474 net1656 n3176 VSS VSS nmos w=1u l=1u
M5475 n3330 net1657 VSS VSS nmos w=1u l=1u
M5476 net1657 n3328 net1658 VSS nmos w=1u l=1u
M5477 net1657 net1655 net1656 VSS nmos w=1u l=1u
M5478 net1658 net1656 VSS VSS nmos w=1u l=1u
M5479 net1657 net1655 net1659 VDD pmos w=2u l=1u
M5480 net1655 n3328 VDD VDD pmos w=2u l=1u
M5481 net1656 n3328 net1657 VDD pmos w=2u l=1u
M5482 net1656 n3176 VDD VDD pmos w=2u l=1u
M5483 n3330 net1657 VDD VDD pmos w=2u l=1u
M5484 net1659 net1656 VDD VDD pmos w=2u l=1u
M5485 n3328 N460 net1660 VSS nmos w=1u l=1u
M5486 net1660 N103 VSS VSS nmos w=1u l=1u
M5487 n3328 N460 VDD VDD pmos w=2u l=1u
M5488 n3328 N103 VDD VDD pmos w=2u l=1u
M5489 n3176 n3175 net1661 VSS nmos w=1u l=1u
M5490 net1661 n3331 VSS VSS nmos w=1u l=1u
M5491 n3176 n3175 VDD VDD pmos w=2u l=1u
M5492 n3176 n3331 VDD VDD pmos w=2u l=1u
M5493 n3175 n3333 net1662 VSS nmos w=1u l=1u
M5494 net1662 n3332 VSS VSS nmos w=1u l=1u
M5495 n3175 n3333 VDD VDD pmos w=2u l=1u
M5496 n3175 n3332 VDD VDD pmos w=2u l=1u
M5497 n3333 n3335 net1663 VSS nmos w=1u l=1u
M5498 net1663 n3334 VSS VSS nmos w=1u l=1u
M5499 n3333 n3335 VDD VDD pmos w=2u l=1u
M5500 n3333 n3334 VDD VDD pmos w=2u l=1u
M5501 n3334 net1664 VSS VSS nmos w=1u l=1u
M5502 net1664 n3336 VSS VSS nmos w=1u l=1u
M5503 net1664 n3337 VSS VSS nmos w=1u l=1u
M5504 net1664 n3337 net1665 VDD pmos w=2u l=1u
M5505 n3334 net1664 VDD VDD pmos w=2u l=1u
M5506 net1665 n3336 VDD VDD pmos w=2u l=1u
M5507 net1666 n3186 VSS VSS nmos w=1u l=1u
M5508 net1667 n3187 VSS VSS nmos w=1u l=1u
M5509 n3332 net1668 VSS VSS nmos w=1u l=1u
M5510 net1668 n3186 net1669 VSS nmos w=1u l=1u
M5511 net1668 net1666 net1667 VSS nmos w=1u l=1u
M5512 net1669 net1667 VSS VSS nmos w=1u l=1u
M5513 net1668 net1666 net1670 VDD pmos w=2u l=1u
M5514 net1666 n3186 VDD VDD pmos w=2u l=1u
M5515 net1667 n3186 net1668 VDD pmos w=2u l=1u
M5516 net1667 n3187 VDD VDD pmos w=2u l=1u
M5517 n3332 net1668 VDD VDD pmos w=2u l=1u
M5518 net1670 net1667 VDD VDD pmos w=2u l=1u
M5519 n3187 n3338 VDD VDD pmos w=2u l=1u
M5520 n3187 n3338 VSS VSS nmos w=1u l=1u
M5521 n3331 n3340 net1671 VSS nmos w=1u l=1u
M5522 net1671 n3339 VSS VSS nmos w=1u l=1u
M5523 n3331 n3340 VDD VDD pmos w=2u l=1u
M5524 n3331 n3339 VDD VDD pmos w=2u l=1u
M5525 net1672 n3338 VSS VSS nmos w=1u l=1u
M5526 net1673 n3186 VSS VSS nmos w=1u l=1u
M5527 n3340 net1674 VSS VSS nmos w=1u l=1u
M5528 net1674 n3338 net1675 VSS nmos w=1u l=1u
M5529 net1674 net1672 net1673 VSS nmos w=1u l=1u
M5530 net1675 net1673 VSS VSS nmos w=1u l=1u
M5531 net1674 net1672 net1676 VDD pmos w=2u l=1u
M5532 net1672 n3338 VDD VDD pmos w=2u l=1u
M5533 net1673 n3338 net1674 VDD pmos w=2u l=1u
M5534 net1673 n3186 VDD VDD pmos w=2u l=1u
M5535 n3340 net1674 VDD VDD pmos w=2u l=1u
M5536 net1676 net1673 VDD VDD pmos w=2u l=1u
M5537 n3338 N443 net1677 VSS nmos w=1u l=1u
M5538 net1677 N120 VSS VSS nmos w=1u l=1u
M5539 n3338 N443 VDD VDD pmos w=2u l=1u
M5540 n3338 N120 VDD VDD pmos w=2u l=1u
M5541 n3186 n3185 net1678 VSS nmos w=1u l=1u
M5542 net1678 n3341 VSS VSS nmos w=1u l=1u
M5543 n3186 n3185 VDD VDD pmos w=2u l=1u
M5544 n3186 n3341 VDD VDD pmos w=2u l=1u
M5545 n3185 n3343 net1679 VSS nmos w=1u l=1u
M5546 net1679 n3342 VSS VSS nmos w=1u l=1u
M5547 n3185 n3343 VDD VDD pmos w=2u l=1u
M5548 n3185 n3342 VDD VDD pmos w=2u l=1u
M5549 n3343 n3345 net1680 VSS nmos w=1u l=1u
M5550 net1680 n3344 VSS VSS nmos w=1u l=1u
M5551 n3343 n3345 VDD VDD pmos w=2u l=1u
M5552 n3343 n3344 VDD VDD pmos w=2u l=1u
M5553 n3344 net1681 VSS VSS nmos w=1u l=1u
M5554 net1681 n3346 VSS VSS nmos w=1u l=1u
M5555 net1681 n3347 VSS VSS nmos w=1u l=1u
M5556 net1681 n3347 net1682 VDD pmos w=2u l=1u
M5557 n3344 net1681 VDD VDD pmos w=2u l=1u
M5558 net1682 n3346 VDD VDD pmos w=2u l=1u
M5559 net1683 n3196 VSS VSS nmos w=1u l=1u
M5560 net1684 n3197 VSS VSS nmos w=1u l=1u
M5561 n3342 net1685 VSS VSS nmos w=1u l=1u
M5562 net1685 n3196 net1686 VSS nmos w=1u l=1u
M5563 net1685 net1683 net1684 VSS nmos w=1u l=1u
M5564 net1686 net1684 VSS VSS nmos w=1u l=1u
M5565 net1685 net1683 net1687 VDD pmos w=2u l=1u
M5566 net1683 n3196 VDD VDD pmos w=2u l=1u
M5567 net1684 n3196 net1685 VDD pmos w=2u l=1u
M5568 net1684 n3197 VDD VDD pmos w=2u l=1u
M5569 n3342 net1685 VDD VDD pmos w=2u l=1u
M5570 net1687 net1684 VDD VDD pmos w=2u l=1u
M5571 n3197 n3348 VDD VDD pmos w=2u l=1u
M5572 n3197 n3348 VSS VSS nmos w=1u l=1u
M5573 n3341 n3350 net1688 VSS nmos w=1u l=1u
M5574 net1688 n3349 VSS VSS nmos w=1u l=1u
M5575 n3341 n3350 VDD VDD pmos w=2u l=1u
M5576 n3341 n3349 VDD VDD pmos w=2u l=1u
M5577 net1689 n3348 VSS VSS nmos w=1u l=1u
M5578 net1690 n3196 VSS VSS nmos w=1u l=1u
M5579 n3350 net1691 VSS VSS nmos w=1u l=1u
M5580 net1691 n3348 net1692 VSS nmos w=1u l=1u
M5581 net1691 net1689 net1690 VSS nmos w=1u l=1u
M5582 net1692 net1690 VSS VSS nmos w=1u l=1u
M5583 net1691 net1689 net1693 VDD pmos w=2u l=1u
M5584 net1689 n3348 VDD VDD pmos w=2u l=1u
M5585 net1690 n3348 net1691 VDD pmos w=2u l=1u
M5586 net1690 n3196 VDD VDD pmos w=2u l=1u
M5587 n3350 net1691 VDD VDD pmos w=2u l=1u
M5588 net1693 net1690 VDD VDD pmos w=2u l=1u
M5589 n3348 N426 net1694 VSS nmos w=1u l=1u
M5590 net1694 N137 VSS VSS nmos w=1u l=1u
M5591 n3348 N426 VDD VDD pmos w=2u l=1u
M5592 n3348 N137 VDD VDD pmos w=2u l=1u
M5593 n3196 n3195 net1695 VSS nmos w=1u l=1u
M5594 net1695 n3351 VSS VSS nmos w=1u l=1u
M5595 n3196 n3195 VDD VDD pmos w=2u l=1u
M5596 n3196 n3351 VDD VDD pmos w=2u l=1u
M5597 n3195 n3353 net1696 VSS nmos w=1u l=1u
M5598 net1696 n3352 VSS VSS nmos w=1u l=1u
M5599 n3195 n3353 VDD VDD pmos w=2u l=1u
M5600 n3195 n3352 VDD VDD pmos w=2u l=1u
M5601 n3353 n3355 net1697 VSS nmos w=1u l=1u
M5602 net1697 n3354 VSS VSS nmos w=1u l=1u
M5603 n3353 n3355 VDD VDD pmos w=2u l=1u
M5604 n3353 n3354 VDD VDD pmos w=2u l=1u
M5605 n3354 net1698 VSS VSS nmos w=1u l=1u
M5606 net1698 n3356 VSS VSS nmos w=1u l=1u
M5607 net1698 n3357 VSS VSS nmos w=1u l=1u
M5608 net1698 n3357 net1699 VDD pmos w=2u l=1u
M5609 n3354 net1698 VDD VDD pmos w=2u l=1u
M5610 net1699 n3356 VDD VDD pmos w=2u l=1u
M5611 net1700 n3206 VSS VSS nmos w=1u l=1u
M5612 net1701 n3207 VSS VSS nmos w=1u l=1u
M5613 n3352 net1702 VSS VSS nmos w=1u l=1u
M5614 net1702 n3206 net1703 VSS nmos w=1u l=1u
M5615 net1702 net1700 net1701 VSS nmos w=1u l=1u
M5616 net1703 net1701 VSS VSS nmos w=1u l=1u
M5617 net1702 net1700 net1704 VDD pmos w=2u l=1u
M5618 net1700 n3206 VDD VDD pmos w=2u l=1u
M5619 net1701 n3206 net1702 VDD pmos w=2u l=1u
M5620 net1701 n3207 VDD VDD pmos w=2u l=1u
M5621 n3352 net1702 VDD VDD pmos w=2u l=1u
M5622 net1704 net1701 VDD VDD pmos w=2u l=1u
M5623 n3207 n3358 VDD VDD pmos w=2u l=1u
M5624 n3207 n3358 VSS VSS nmos w=1u l=1u
M5625 n3351 n3360 net1705 VSS nmos w=1u l=1u
M5626 net1705 n3359 VSS VSS nmos w=1u l=1u
M5627 n3351 n3360 VDD VDD pmos w=2u l=1u
M5628 n3351 n3359 VDD VDD pmos w=2u l=1u
M5629 net1706 n3358 VSS VSS nmos w=1u l=1u
M5630 net1707 n3206 VSS VSS nmos w=1u l=1u
M5631 n3360 net1708 VSS VSS nmos w=1u l=1u
M5632 net1708 n3358 net1709 VSS nmos w=1u l=1u
M5633 net1708 net1706 net1707 VSS nmos w=1u l=1u
M5634 net1709 net1707 VSS VSS nmos w=1u l=1u
M5635 net1708 net1706 net1710 VDD pmos w=2u l=1u
M5636 net1706 n3358 VDD VDD pmos w=2u l=1u
M5637 net1707 n3358 net1708 VDD pmos w=2u l=1u
M5638 net1707 n3206 VDD VDD pmos w=2u l=1u
M5639 n3360 net1708 VDD VDD pmos w=2u l=1u
M5640 net1710 net1707 VDD VDD pmos w=2u l=1u
M5641 n3358 N409 net1711 VSS nmos w=1u l=1u
M5642 net1711 N154 VSS VSS nmos w=1u l=1u
M5643 n3358 N409 VDD VDD pmos w=2u l=1u
M5644 n3358 N154 VDD VDD pmos w=2u l=1u
M5645 n3206 n3205 net1712 VSS nmos w=1u l=1u
M5646 net1712 n3361 VSS VSS nmos w=1u l=1u
M5647 n3206 n3205 VDD VDD pmos w=2u l=1u
M5648 n3206 n3361 VDD VDD pmos w=2u l=1u
M5649 n3205 n3363 net1713 VSS nmos w=1u l=1u
M5650 net1713 n3362 VSS VSS nmos w=1u l=1u
M5651 n3205 n3363 VDD VDD pmos w=2u l=1u
M5652 n3205 n3362 VDD VDD pmos w=2u l=1u
M5653 n3363 n3365 net1714 VSS nmos w=1u l=1u
M5654 net1714 n3364 VSS VSS nmos w=1u l=1u
M5655 n3363 n3365 VDD VDD pmos w=2u l=1u
M5656 n3363 n3364 VDD VDD pmos w=2u l=1u
M5657 n3364 net1715 VSS VSS nmos w=1u l=1u
M5658 net1715 n3366 VSS VSS nmos w=1u l=1u
M5659 net1715 n3367 VSS VSS nmos w=1u l=1u
M5660 net1715 n3367 net1716 VDD pmos w=2u l=1u
M5661 n3364 net1715 VDD VDD pmos w=2u l=1u
M5662 net1716 n3366 VDD VDD pmos w=2u l=1u
M5663 net1717 n3216 VSS VSS nmos w=1u l=1u
M5664 net1718 n3217 VSS VSS nmos w=1u l=1u
M5665 n3362 net1719 VSS VSS nmos w=1u l=1u
M5666 net1719 n3216 net1720 VSS nmos w=1u l=1u
M5667 net1719 net1717 net1718 VSS nmos w=1u l=1u
M5668 net1720 net1718 VSS VSS nmos w=1u l=1u
M5669 net1719 net1717 net1721 VDD pmos w=2u l=1u
M5670 net1717 n3216 VDD VDD pmos w=2u l=1u
M5671 net1718 n3216 net1719 VDD pmos w=2u l=1u
M5672 net1718 n3217 VDD VDD pmos w=2u l=1u
M5673 n3362 net1719 VDD VDD pmos w=2u l=1u
M5674 net1721 net1718 VDD VDD pmos w=2u l=1u
M5675 n3217 n3368 VDD VDD pmos w=2u l=1u
M5676 n3217 n3368 VSS VSS nmos w=1u l=1u
M5677 n3361 n3370 net1722 VSS nmos w=1u l=1u
M5678 net1722 n3369 VSS VSS nmos w=1u l=1u
M5679 n3361 n3370 VDD VDD pmos w=2u l=1u
M5680 n3361 n3369 VDD VDD pmos w=2u l=1u
M5681 net1723 n3368 VSS VSS nmos w=1u l=1u
M5682 net1724 n3216 VSS VSS nmos w=1u l=1u
M5683 n3370 net1725 VSS VSS nmos w=1u l=1u
M5684 net1725 n3368 net1726 VSS nmos w=1u l=1u
M5685 net1725 net1723 net1724 VSS nmos w=1u l=1u
M5686 net1726 net1724 VSS VSS nmos w=1u l=1u
M5687 net1725 net1723 net1727 VDD pmos w=2u l=1u
M5688 net1723 n3368 VDD VDD pmos w=2u l=1u
M5689 net1724 n3368 net1725 VDD pmos w=2u l=1u
M5690 net1724 n3216 VDD VDD pmos w=2u l=1u
M5691 n3370 net1725 VDD VDD pmos w=2u l=1u
M5692 net1727 net1724 VDD VDD pmos w=2u l=1u
M5693 n3368 N392 net1728 VSS nmos w=1u l=1u
M5694 net1728 N171 VSS VSS nmos w=1u l=1u
M5695 n3368 N392 VDD VDD pmos w=2u l=1u
M5696 n3368 N171 VDD VDD pmos w=2u l=1u
M5697 n3216 n3215 net1729 VSS nmos w=1u l=1u
M5698 net1729 n3371 VSS VSS nmos w=1u l=1u
M5699 n3216 n3215 VDD VDD pmos w=2u l=1u
M5700 n3216 n3371 VDD VDD pmos w=2u l=1u
M5701 n3215 n3373 net1730 VSS nmos w=1u l=1u
M5702 net1730 n3372 VSS VSS nmos w=1u l=1u
M5703 n3215 n3373 VDD VDD pmos w=2u l=1u
M5704 n3215 n3372 VDD VDD pmos w=2u l=1u
M5705 n3373 n3375 net1731 VSS nmos w=1u l=1u
M5706 net1731 n3374 VSS VSS nmos w=1u l=1u
M5707 n3373 n3375 VDD VDD pmos w=2u l=1u
M5708 n3373 n3374 VDD VDD pmos w=2u l=1u
M5709 n3374 n3377 net1732 VSS nmos w=1u l=1u
M5710 net1732 n3376 VSS VSS nmos w=1u l=1u
M5711 n3374 n3377 VDD VDD pmos w=2u l=1u
M5712 n3374 n3376 VDD VDD pmos w=2u l=1u
M5713 net1733 n3226 VSS VSS nmos w=1u l=1u
M5714 net1734 n3227 VSS VSS nmos w=1u l=1u
M5715 n3372 net1735 VSS VSS nmos w=1u l=1u
M5716 net1735 n3226 net1736 VSS nmos w=1u l=1u
M5717 net1735 net1733 net1734 VSS nmos w=1u l=1u
M5718 net1736 net1734 VSS VSS nmos w=1u l=1u
M5719 net1735 net1733 net1737 VDD pmos w=2u l=1u
M5720 net1733 n3226 VDD VDD pmos w=2u l=1u
M5721 net1734 n3226 net1735 VDD pmos w=2u l=1u
M5722 net1734 n3227 VDD VDD pmos w=2u l=1u
M5723 n3372 net1735 VDD VDD pmos w=2u l=1u
M5724 net1737 net1734 VDD VDD pmos w=2u l=1u
M5725 n3227 n3378 VDD VDD pmos w=2u l=1u
M5726 n3227 n3378 VSS VSS nmos w=1u l=1u
M5727 n3371 n3380 net1738 VSS nmos w=1u l=1u
M5728 net1738 n3379 VSS VSS nmos w=1u l=1u
M5729 n3371 n3380 VDD VDD pmos w=2u l=1u
M5730 n3371 n3379 VDD VDD pmos w=2u l=1u
M5731 net1739 n3378 VSS VSS nmos w=1u l=1u
M5732 net1740 n3226 VSS VSS nmos w=1u l=1u
M5733 n3380 net1741 VSS VSS nmos w=1u l=1u
M5734 net1741 n3378 net1742 VSS nmos w=1u l=1u
M5735 net1741 net1739 net1740 VSS nmos w=1u l=1u
M5736 net1742 net1740 VSS VSS nmos w=1u l=1u
M5737 net1741 net1739 net1743 VDD pmos w=2u l=1u
M5738 net1739 n3378 VDD VDD pmos w=2u l=1u
M5739 net1740 n3378 net1741 VDD pmos w=2u l=1u
M5740 net1740 n3226 VDD VDD pmos w=2u l=1u
M5741 n3380 net1741 VDD VDD pmos w=2u l=1u
M5742 net1743 net1740 VDD VDD pmos w=2u l=1u
M5743 n3378 N375 net1744 VSS nmos w=1u l=1u
M5744 net1744 N188 VSS VSS nmos w=1u l=1u
M5745 n3378 N375 VDD VDD pmos w=2u l=1u
M5746 n3378 N188 VDD VDD pmos w=2u l=1u
M5747 n3226 n3225 net1745 VSS nmos w=1u l=1u
M5748 net1745 n3381 VSS VSS nmos w=1u l=1u
M5749 n3226 n3225 VDD VDD pmos w=2u l=1u
M5750 n3226 n3381 VDD VDD pmos w=2u l=1u
M5751 n3225 n3383 net1746 VSS nmos w=1u l=1u
M5752 net1746 n3382 VSS VSS nmos w=1u l=1u
M5753 n3225 n3383 VDD VDD pmos w=2u l=1u
M5754 n3225 n3382 VDD VDD pmos w=2u l=1u
M5755 n3383 n3385 net1747 VSS nmos w=1u l=1u
M5756 net1747 n3384 VSS VSS nmos w=1u l=1u
M5757 n3383 n3385 VDD VDD pmos w=2u l=1u
M5758 n3383 n3384 VDD VDD pmos w=2u l=1u
M5759 n3384 net1748 VSS VSS nmos w=1u l=1u
M5760 net1748 n3386 VSS VSS nmos w=1u l=1u
M5761 net1748 n3387 VSS VSS nmos w=1u l=1u
M5762 net1748 n3387 net1749 VDD pmos w=2u l=1u
M5763 n3384 net1748 VDD VDD pmos w=2u l=1u
M5764 net1749 n3386 VDD VDD pmos w=2u l=1u
M5765 net1750 n3236 VSS VSS nmos w=1u l=1u
M5766 net1751 n3237 VSS VSS nmos w=1u l=1u
M5767 n3382 net1752 VSS VSS nmos w=1u l=1u
M5768 net1752 n3236 net1753 VSS nmos w=1u l=1u
M5769 net1752 net1750 net1751 VSS nmos w=1u l=1u
M5770 net1753 net1751 VSS VSS nmos w=1u l=1u
M5771 net1752 net1750 net1754 VDD pmos w=2u l=1u
M5772 net1750 n3236 VDD VDD pmos w=2u l=1u
M5773 net1751 n3236 net1752 VDD pmos w=2u l=1u
M5774 net1751 n3237 VDD VDD pmos w=2u l=1u
M5775 n3382 net1752 VDD VDD pmos w=2u l=1u
M5776 net1754 net1751 VDD VDD pmos w=2u l=1u
M5777 n3237 n3388 VDD VDD pmos w=2u l=1u
M5778 n3237 n3388 VSS VSS nmos w=1u l=1u
M5779 n3381 n3390 net1755 VSS nmos w=1u l=1u
M5780 net1755 n3389 VSS VSS nmos w=1u l=1u
M5781 n3381 n3390 VDD VDD pmos w=2u l=1u
M5782 n3381 n3389 VDD VDD pmos w=2u l=1u
M5783 net1756 n3388 VSS VSS nmos w=1u l=1u
M5784 net1757 n3236 VSS VSS nmos w=1u l=1u
M5785 n3390 net1758 VSS VSS nmos w=1u l=1u
M5786 net1758 n3388 net1759 VSS nmos w=1u l=1u
M5787 net1758 net1756 net1757 VSS nmos w=1u l=1u
M5788 net1759 net1757 VSS VSS nmos w=1u l=1u
M5789 net1758 net1756 net1760 VDD pmos w=2u l=1u
M5790 net1756 n3388 VDD VDD pmos w=2u l=1u
M5791 net1757 n3388 net1758 VDD pmos w=2u l=1u
M5792 net1757 n3236 VDD VDD pmos w=2u l=1u
M5793 n3390 net1758 VDD VDD pmos w=2u l=1u
M5794 net1760 net1757 VDD VDD pmos w=2u l=1u
M5795 n3388 N358 net1761 VSS nmos w=1u l=1u
M5796 net1761 N205 VSS VSS nmos w=1u l=1u
M5797 n3388 N358 VDD VDD pmos w=2u l=1u
M5798 n3388 N205 VDD VDD pmos w=2u l=1u
M5799 n3236 n3235 net1762 VSS nmos w=1u l=1u
M5800 net1762 n3391 VSS VSS nmos w=1u l=1u
M5801 n3236 n3235 VDD VDD pmos w=2u l=1u
M5802 n3236 n3391 VDD VDD pmos w=2u l=1u
M5803 n3235 n3393 net1763 VSS nmos w=1u l=1u
M5804 net1763 n3392 VSS VSS nmos w=1u l=1u
M5805 n3235 n3393 VDD VDD pmos w=2u l=1u
M5806 n3235 n3392 VDD VDD pmos w=2u l=1u
M5807 n3393 n3395 net1764 VSS nmos w=1u l=1u
M5808 net1764 n3394 VSS VSS nmos w=1u l=1u
M5809 n3393 n3395 VDD VDD pmos w=2u l=1u
M5810 n3393 n3394 VDD VDD pmos w=2u l=1u
M5811 n3394 net1765 VSS VSS nmos w=1u l=1u
M5812 net1765 n3396 VSS VSS nmos w=1u l=1u
M5813 net1765 n3397 VSS VSS nmos w=1u l=1u
M5814 net1765 n3397 net1766 VDD pmos w=2u l=1u
M5815 n3394 net1765 VDD VDD pmos w=2u l=1u
M5816 net1766 n3396 VDD VDD pmos w=2u l=1u
M5817 net1767 n3247 VSS VSS nmos w=1u l=1u
M5818 net1768 n3248 VSS VSS nmos w=1u l=1u
M5819 n3392 net1769 VSS VSS nmos w=1u l=1u
M5820 net1769 n3247 net1770 VSS nmos w=1u l=1u
M5821 net1769 net1767 net1768 VSS nmos w=1u l=1u
M5822 net1770 net1768 VSS VSS nmos w=1u l=1u
M5823 net1769 net1767 net1771 VDD pmos w=2u l=1u
M5824 net1767 n3247 VDD VDD pmos w=2u l=1u
M5825 net1768 n3247 net1769 VDD pmos w=2u l=1u
M5826 net1768 n3248 VDD VDD pmos w=2u l=1u
M5827 n3392 net1769 VDD VDD pmos w=2u l=1u
M5828 net1771 net1768 VDD VDD pmos w=2u l=1u
M5829 n3247 n3398 VDD VDD pmos w=2u l=1u
M5830 n3247 n3398 VSS VSS nmos w=1u l=1u
M5831 n3391 n3400 net1772 VSS nmos w=1u l=1u
M5832 net1772 n3399 VSS VSS nmos w=1u l=1u
M5833 n3391 n3400 VDD VDD pmos w=2u l=1u
M5834 n3391 n3399 VDD VDD pmos w=2u l=1u
M5835 net1773 n3248 VSS VSS nmos w=1u l=1u
M5836 net1774 n3398 VSS VSS nmos w=1u l=1u
M5837 n3400 net1775 VSS VSS nmos w=1u l=1u
M5838 net1775 n3248 net1776 VSS nmos w=1u l=1u
M5839 net1775 net1773 net1774 VSS nmos w=1u l=1u
M5840 net1776 net1774 VSS VSS nmos w=1u l=1u
M5841 net1775 net1773 net1777 VDD pmos w=2u l=1u
M5842 net1773 n3248 VDD VDD pmos w=2u l=1u
M5843 net1774 n3248 net1775 VDD pmos w=2u l=1u
M5844 net1774 n3398 VDD VDD pmos w=2u l=1u
M5845 n3400 net1775 VDD VDD pmos w=2u l=1u
M5846 net1777 net1774 VDD VDD pmos w=2u l=1u
M5847 n3248 N341 net1778 VSS nmos w=1u l=1u
M5848 net1778 N222 VSS VSS nmos w=1u l=1u
M5849 n3248 N341 VDD VDD pmos w=2u l=1u
M5850 n3248 N222 VDD VDD pmos w=2u l=1u
M5851 n3398 n3245 net1779 VSS nmos w=1u l=1u
M5852 net1779 n3401 VSS VSS nmos w=1u l=1u
M5853 n3398 n3245 VDD VDD pmos w=2u l=1u
M5854 n3398 n3401 VDD VDD pmos w=2u l=1u
M5855 n3245 n3249 VDD VDD pmos w=2u l=1u
M5856 n3245 n3249 VSS VSS nmos w=1u l=1u
M5857 n3249 n3403 VSS VSS nmos w=1u l=1u
M5858 n3249 n3402 VSS VSS nmos w=1u l=1u
M5859 n3249 n3403 net1780 VDD pmos w=2u l=1u
M5860 net1780 n3402 VDD VDD pmos w=2u l=1u
M5861 n3401 n3402 net1781 VSS nmos w=1u l=1u
M5862 net1781 n3403 VSS VSS nmos w=1u l=1u
M5863 n3401 n3402 VDD VDD pmos w=2u l=1u
M5864 n3401 n3403 VDD VDD pmos w=2u l=1u
M5865 n3402 n3404 net1782 VSS nmos w=1u l=1u
M5866 net1782 n3260 VSS VSS nmos w=1u l=1u
M5867 n3402 n3404 VDD VDD pmos w=2u l=1u
M5868 n3402 n3260 VDD VDD pmos w=2u l=1u
M5869 n3404 N324 net1783 VSS nmos w=1u l=1u
M5870 net1783 n3405 VSS VSS nmos w=1u l=1u
M5871 n3404 N324 VDD VDD pmos w=2u l=1u
M5872 n3404 n3405 VDD VDD pmos w=2u l=1u
M5873 n3405 n3407 VSS VSS nmos w=1u l=1u
M5874 n3405 n3406 VSS VSS nmos w=1u l=1u
M5875 n3405 n3407 net1784 VDD pmos w=2u l=1u
M5876 net1784 n3406 VDD VDD pmos w=2u l=1u
M5877 n3407 n3409 VSS VSS nmos w=1u l=1u
M5878 n3407 n3408 VSS VSS nmos w=1u l=1u
M5879 n3407 n3409 net1785 VDD pmos w=2u l=1u
M5880 net1785 n3408 VDD VDD pmos w=2u l=1u
M5881 n3409 n2270 net1786 VSS nmos w=1u l=1u
M5882 net1786 n3410 VSS VSS nmos w=1u l=1u
M5883 n3409 n2270 VDD VDD pmos w=2u l=1u
M5884 n3409 n3410 VDD VDD pmos w=2u l=1u
M5885 n3410 n3411 net1787 VSS nmos w=1u l=1u
M5886 net1787 N239 VSS VSS nmos w=1u l=1u
M5887 n3410 n3411 VDD VDD pmos w=2u l=1u
M5888 n3410 N239 VDD VDD pmos w=2u l=1u
M5889 n3408 n3263 VDD VDD pmos w=2u l=1u
M5890 n3408 n3263 VSS VSS nmos w=1u l=1u
M5891 n3406 n3263 VSS VSS nmos w=1u l=1u
M5892 n3406 N307 VSS VSS nmos w=1u l=1u
M5893 n3406 n3263 net1788 VDD pmos w=2u l=1u
M5894 net1788 N307 VDD VDD pmos w=2u l=1u
M5895 n3260 n3413 net1789 VSS nmos w=1u l=1u
M5896 net1789 n3412 VSS VSS nmos w=1u l=1u
M5897 n3260 n3413 VDD VDD pmos w=2u l=1u
M5898 n3260 n3412 VDD VDD pmos w=2u l=1u
M5899 n3413 N239 net1790 VSS nmos w=1u l=1u
M5900 net1790 N324 VSS VSS nmos w=1u l=1u
M5901 n3413 N239 VDD VDD pmos w=2u l=1u
M5902 n3413 N324 VDD VDD pmos w=2u l=1u
M5903 net1791 n3262 VSS VSS nmos w=1u l=1u
M5904 net1792 n3263 VSS VSS nmos w=1u l=1u
M5905 n3412 net1793 VSS VSS nmos w=1u l=1u
M5906 net1793 n3262 net1794 VSS nmos w=1u l=1u
M5907 net1793 net1791 net1792 VSS nmos w=1u l=1u
M5908 net1794 net1792 VSS VSS nmos w=1u l=1u
M5909 net1793 net1791 net1795 VDD pmos w=2u l=1u
M5910 net1791 n3262 VDD VDD pmos w=2u l=1u
M5911 net1792 n3262 net1793 VDD pmos w=2u l=1u
M5912 net1792 n3263 VDD VDD pmos w=2u l=1u
M5913 n3412 net1793 VDD VDD pmos w=2u l=1u
M5914 net1795 net1792 VDD VDD pmos w=2u l=1u
M5915 n3262 N256 net1796 VSS nmos w=1u l=1u
M5916 net1796 N307 VSS VSS nmos w=1u l=1u
M5917 n3262 N256 VDD VDD pmos w=2u l=1u
M5918 n3262 N307 VDD VDD pmos w=2u l=1u
M5919 n3263 N290 net1797 VSS nmos w=1u l=1u
M5920 net1797 n3414 VSS VSS nmos w=1u l=1u
M5921 n3263 N290 VDD VDD pmos w=2u l=1u
M5922 n3263 n3414 VDD VDD pmos w=2u l=1u
M5923 n3414 net1798 VSS VSS nmos w=1u l=1u
M5924 net1799 N256 VSS VSS nmos w=1u l=1u
M5925 net1798 n3415 net1799 VSS nmos w=1u l=1u
M5926 net1798 N256 VDD VDD pmos w=2u l=1u
M5927 net1798 n3415 VDD VDD pmos w=2u l=1u
M5928 n3414 net1798 VDD VDD pmos w=2u l=1u
M5929 n3403 n3417 VSS VSS nmos w=1u l=1u
M5930 n3403 n3416 VSS VSS nmos w=1u l=1u
M5931 n3403 n3417 net1800 VDD pmos w=2u l=1u
M5932 net1800 n3416 VDD VDD pmos w=2u l=1u
M5933 n3417 n3418 VDD VDD pmos w=2u l=1u
M5934 n3417 n3418 VSS VSS nmos w=1u l=1u
M5935 n3399 n3420 VSS VSS nmos w=1u l=1u
M5936 n3399 n3419 VSS VSS nmos w=1u l=1u
M5937 n3399 n3420 net1801 VDD pmos w=2u l=1u
M5938 net1801 n3419 VDD VDD pmos w=2u l=1u
M5939 n3420 n3396 VSS VSS nmos w=1u l=1u
M5940 n3420 n3397 VSS VSS nmos w=1u l=1u
M5941 n3420 n3396 net1802 VDD pmos w=2u l=1u
M5942 net1802 n3397 VDD VDD pmos w=2u l=1u
M5943 n3419 n3395 VDD VDD pmos w=2u l=1u
M5944 n3419 n3395 VSS VSS nmos w=1u l=1u
M5945 n3389 n3422 VSS VSS nmos w=1u l=1u
M5946 n3389 n3421 VSS VSS nmos w=1u l=1u
M5947 n3389 n3422 net1803 VDD pmos w=2u l=1u
M5948 net1803 n3421 VDD VDD pmos w=2u l=1u
M5949 n3422 n3386 VSS VSS nmos w=1u l=1u
M5950 n3422 n3387 VSS VSS nmos w=1u l=1u
M5951 n3422 n3386 net1804 VDD pmos w=2u l=1u
M5952 net1804 n3387 VDD VDD pmos w=2u l=1u
M5953 n3421 n3385 VDD VDD pmos w=2u l=1u
M5954 n3421 n3385 VSS VSS nmos w=1u l=1u
M5955 n3379 n3424 VSS VSS nmos w=1u l=1u
M5956 n3379 n3423 VSS VSS nmos w=1u l=1u
M5957 n3379 n3424 net1805 VDD pmos w=2u l=1u
M5958 net1805 n3423 VDD VDD pmos w=2u l=1u
M5959 n3424 net1806 VSS VSS nmos w=1u l=1u
M5960 net1807 n3376 VSS VSS nmos w=1u l=1u
M5961 net1806 n3377 net1807 VSS nmos w=1u l=1u
M5962 net1806 n3376 VDD VDD pmos w=2u l=1u
M5963 net1806 n3377 VDD VDD pmos w=2u l=1u
M5964 n3424 net1806 VDD VDD pmos w=2u l=1u
M5965 n3423 n3375 VDD VDD pmos w=2u l=1u
M5966 n3423 n3375 VSS VSS nmos w=1u l=1u
M5967 n3369 n3426 VSS VSS nmos w=1u l=1u
M5968 n3369 n3425 VSS VSS nmos w=1u l=1u
M5969 n3369 n3426 net1808 VDD pmos w=2u l=1u
M5970 net1808 n3425 VDD VDD pmos w=2u l=1u
M5971 n3426 n3366 VSS VSS nmos w=1u l=1u
M5972 n3426 n3367 VSS VSS nmos w=1u l=1u
M5973 n3426 n3366 net1809 VDD pmos w=2u l=1u
M5974 net1809 n3367 VDD VDD pmos w=2u l=1u
M5975 n3425 n3365 VDD VDD pmos w=2u l=1u
M5976 n3425 n3365 VSS VSS nmos w=1u l=1u
M5977 n3359 n3428 VSS VSS nmos w=1u l=1u
M5978 n3359 n3427 VSS VSS nmos w=1u l=1u
M5979 n3359 n3428 net1810 VDD pmos w=2u l=1u
M5980 net1810 n3427 VDD VDD pmos w=2u l=1u
M5981 n3428 n3356 VSS VSS nmos w=1u l=1u
M5982 n3428 n3357 VSS VSS nmos w=1u l=1u
M5983 n3428 n3356 net1811 VDD pmos w=2u l=1u
M5984 net1811 n3357 VDD VDD pmos w=2u l=1u
M5985 n3427 n3355 VDD VDD pmos w=2u l=1u
M5986 n3427 n3355 VSS VSS nmos w=1u l=1u
M5987 n3349 n3430 VSS VSS nmos w=1u l=1u
M5988 n3349 n3429 VSS VSS nmos w=1u l=1u
M5989 n3349 n3430 net1812 VDD pmos w=2u l=1u
M5990 net1812 n3429 VDD VDD pmos w=2u l=1u
M5991 n3430 n3346 VSS VSS nmos w=1u l=1u
M5992 n3430 n3347 VSS VSS nmos w=1u l=1u
M5993 n3430 n3346 net1813 VDD pmos w=2u l=1u
M5994 net1813 n3347 VDD VDD pmos w=2u l=1u
M5995 n3429 n3345 VDD VDD pmos w=2u l=1u
M5996 n3429 n3345 VSS VSS nmos w=1u l=1u
M5997 n3339 n3432 VSS VSS nmos w=1u l=1u
M5998 n3339 n3431 VSS VSS nmos w=1u l=1u
M5999 n3339 n3432 net1814 VDD pmos w=2u l=1u
M6000 net1814 n3431 VDD VDD pmos w=2u l=1u
M6001 n3432 n3336 VSS VSS nmos w=1u l=1u
M6002 n3432 n3337 VSS VSS nmos w=1u l=1u
M6003 n3432 n3336 net1815 VDD pmos w=2u l=1u
M6004 net1815 n3337 VDD VDD pmos w=2u l=1u
M6005 n3431 n3335 VDD VDD pmos w=2u l=1u
M6006 n3431 n3335 VSS VSS nmos w=1u l=1u
M6007 n3329 n3434 VSS VSS nmos w=1u l=1u
M6008 n3329 n3433 VSS VSS nmos w=1u l=1u
M6009 n3329 n3434 net1816 VDD pmos w=2u l=1u
M6010 net1816 n3433 VDD VDD pmos w=2u l=1u
M6011 n3434 n3326 VSS VSS nmos w=1u l=1u
M6012 n3434 n3327 VSS VSS nmos w=1u l=1u
M6013 n3434 n3326 net1817 VDD pmos w=2u l=1u
M6014 net1817 n3327 VDD VDD pmos w=2u l=1u
M6015 n3433 n3325 VDD VDD pmos w=2u l=1u
M6016 n3433 n3325 VSS VSS nmos w=1u l=1u
M6017 n3319 n3436 VSS VSS nmos w=1u l=1u
M6018 n3319 n3435 VSS VSS nmos w=1u l=1u
M6019 n3319 n3436 net1818 VDD pmos w=2u l=1u
M6020 net1818 n3435 VDD VDD pmos w=2u l=1u
M6021 n3436 n3316 VSS VSS nmos w=1u l=1u
M6022 n3436 n3317 VSS VSS nmos w=1u l=1u
M6023 n3436 n3316 net1819 VDD pmos w=2u l=1u
M6024 net1819 n3317 VDD VDD pmos w=2u l=1u
M6025 n3435 n3315 VDD VDD pmos w=2u l=1u
M6026 n3435 n3315 VSS VSS nmos w=1u l=1u
M6027 n3309 n3438 VSS VSS nmos w=1u l=1u
M6028 n3309 n3437 VSS VSS nmos w=1u l=1u
M6029 n3309 n3438 net1820 VDD pmos w=2u l=1u
M6030 net1820 n3437 VDD VDD pmos w=2u l=1u
M6031 n3438 n3306 VSS VSS nmos w=1u l=1u
M6032 n3438 n3307 VSS VSS nmos w=1u l=1u
M6033 n3438 n3306 net1821 VDD pmos w=2u l=1u
M6034 net1821 n3307 VDD VDD pmos w=2u l=1u
M6035 n3437 n3305 VDD VDD pmos w=2u l=1u
M6036 n3437 n3305 VSS VSS nmos w=1u l=1u
M6037 n3299 n3440 VSS VSS nmos w=1u l=1u
M6038 n3299 n3439 VSS VSS nmos w=1u l=1u
M6039 n3299 n3440 net1822 VDD pmos w=2u l=1u
M6040 net1822 n3439 VDD VDD pmos w=2u l=1u
M6041 n3440 n3296 VSS VSS nmos w=1u l=1u
M6042 n3440 n3297 VSS VSS nmos w=1u l=1u
M6043 n3440 n3296 net1823 VDD pmos w=2u l=1u
M6044 net1823 n3297 VDD VDD pmos w=2u l=1u
M6045 n3439 n3295 VDD VDD pmos w=2u l=1u
M6046 n3439 n3295 VSS VSS nmos w=1u l=1u
M6047 n3140 N528 net1824 VSS nmos w=1u l=1u
M6048 net1824 N35 VSS VSS nmos w=1u l=1u
M6049 n3140 N528 VDD VDD pmos w=2u l=1u
M6050 n3140 N35 VDD VDD pmos w=2u l=1u
M6051 N6150 n3442 VSS VSS nmos w=1u l=1u
M6052 N6150 n3441 VSS VSS nmos w=1u l=1u
M6053 N6150 n3442 net1825 VDD pmos w=2u l=1u
M6054 net1825 n3441 VDD VDD pmos w=2u l=1u
M6055 n3442 n3444 VSS VSS nmos w=1u l=1u
M6056 n3442 n3443 VSS VSS nmos w=1u l=1u
M6057 n3442 n3444 net1826 VDD pmos w=2u l=1u
M6058 net1826 n3443 VDD VDD pmos w=2u l=1u
M6059 n3441 n3286 VDD VDD pmos w=2u l=1u
M6060 n3441 n3286 VSS VSS nmos w=1u l=1u
M6061 n3286 n3444 net1827 VSS nmos w=1u l=1u
M6062 net1827 n3443 VSS VSS nmos w=1u l=1u
M6063 n3286 n3444 VDD VDD pmos w=2u l=1u
M6064 n3286 n3443 VDD VDD pmos w=2u l=1u
M6065 net1828 n3289 VSS VSS nmos w=1u l=1u
M6066 net1829 n3445 VSS VSS nmos w=1u l=1u
M6067 n3444 net1830 VSS VSS nmos w=1u l=1u
M6068 net1830 n3289 net1831 VSS nmos w=1u l=1u
M6069 net1830 net1828 net1829 VSS nmos w=1u l=1u
M6070 net1831 net1829 VSS VSS nmos w=1u l=1u
M6071 net1830 net1828 net1832 VDD pmos w=2u l=1u
M6072 net1828 n3289 VDD VDD pmos w=2u l=1u
M6073 net1829 n3289 net1830 VDD pmos w=2u l=1u
M6074 net1829 n3445 VDD VDD pmos w=2u l=1u
M6075 n3444 net1830 VDD VDD pmos w=2u l=1u
M6076 net1832 net1829 VDD VDD pmos w=2u l=1u
M6077 n3289 net1833 VSS VSS nmos w=1u l=1u
M6078 net1834 n3288 VSS VSS nmos w=1u l=1u
M6079 net1833 n3446 net1834 VSS nmos w=1u l=1u
M6080 net1833 n3288 VDD VDD pmos w=2u l=1u
M6081 net1833 n3446 VDD VDD pmos w=2u l=1u
M6082 n3289 net1833 VDD VDD pmos w=2u l=1u
M6083 n3288 n3448 net1835 VSS nmos w=1u l=1u
M6084 net1835 n3447 VSS VSS nmos w=1u l=1u
M6085 n3288 n3448 VDD VDD pmos w=2u l=1u
M6086 n3288 n3447 VDD VDD pmos w=2u l=1u
M6087 n3448 n3450 net1836 VSS nmos w=1u l=1u
M6088 net1836 n3449 VSS VSS nmos w=1u l=1u
M6089 n3448 n3450 VDD VDD pmos w=2u l=1u
M6090 n3448 n3449 VDD VDD pmos w=2u l=1u
M6091 n3449 net1837 VSS VSS nmos w=1u l=1u
M6092 net1837 n3451 VSS VSS nmos w=1u l=1u
M6093 net1837 n3452 VSS VSS nmos w=1u l=1u
M6094 net1837 n3452 net1838 VDD pmos w=2u l=1u
M6095 n3449 net1837 VDD VDD pmos w=2u l=1u
M6096 net1838 n3451 VDD VDD pmos w=2u l=1u
M6097 net1839 n3296 VSS VSS nmos w=1u l=1u
M6098 net1840 n3297 VSS VSS nmos w=1u l=1u
M6099 n3447 net1841 VSS VSS nmos w=1u l=1u
M6100 net1841 n3296 net1842 VSS nmos w=1u l=1u
M6101 net1841 net1839 net1840 VSS nmos w=1u l=1u
M6102 net1842 net1840 VSS VSS nmos w=1u l=1u
M6103 net1841 net1839 net1843 VDD pmos w=2u l=1u
M6104 net1839 n3296 VDD VDD pmos w=2u l=1u
M6105 net1840 n3296 net1841 VDD pmos w=2u l=1u
M6106 net1840 n3297 VDD VDD pmos w=2u l=1u
M6107 n3447 net1841 VDD VDD pmos w=2u l=1u
M6108 net1843 net1840 VDD VDD pmos w=2u l=1u
M6109 n3446 n3454 net1844 VSS nmos w=1u l=1u
M6110 net1844 n3453 VSS VSS nmos w=1u l=1u
M6111 n3446 n3454 VDD VDD pmos w=2u l=1u
M6112 n3446 n3453 VDD VDD pmos w=2u l=1u
M6113 net1845 n3297 VSS VSS nmos w=1u l=1u
M6114 net1846 n3455 VSS VSS nmos w=1u l=1u
M6115 n3454 net1847 VSS VSS nmos w=1u l=1u
M6116 net1847 n3297 net1848 VSS nmos w=1u l=1u
M6117 net1847 net1845 net1846 VSS nmos w=1u l=1u
M6118 net1848 net1846 VSS VSS nmos w=1u l=1u
M6119 net1847 net1845 net1849 VDD pmos w=2u l=1u
M6120 net1845 n3297 VDD VDD pmos w=2u l=1u
M6121 net1846 n3297 net1847 VDD pmos w=2u l=1u
M6122 net1846 n3455 VDD VDD pmos w=2u l=1u
M6123 n3454 net1847 VDD VDD pmos w=2u l=1u
M6124 net1849 net1846 VDD VDD pmos w=2u l=1u
M6125 n3297 n2232 VSS VSS nmos w=1u l=1u
M6126 n3297 n3456 VSS VSS nmos w=1u l=1u
M6127 n3297 n2232 net1850 VDD pmos w=2u l=1u
M6128 net1850 n3456 VDD VDD pmos w=2u l=1u
M6129 n3455 n3296 VDD VDD pmos w=2u l=1u
M6130 n3455 n3296 VSS VSS nmos w=1u l=1u
M6131 n3296 n3295 net1851 VSS nmos w=1u l=1u
M6132 net1851 n3457 VSS VSS nmos w=1u l=1u
M6133 n3296 n3295 VDD VDD pmos w=2u l=1u
M6134 n3296 n3457 VDD VDD pmos w=2u l=1u
M6135 n3295 n3459 net1852 VSS nmos w=1u l=1u
M6136 net1852 n3458 VSS VSS nmos w=1u l=1u
M6137 n3295 n3459 VDD VDD pmos w=2u l=1u
M6138 n3295 n3458 VDD VDD pmos w=2u l=1u
M6139 n3459 n3461 net1853 VSS nmos w=1u l=1u
M6140 net1853 n3460 VSS VSS nmos w=1u l=1u
M6141 n3459 n3461 VDD VDD pmos w=2u l=1u
M6142 n3459 n3460 VDD VDD pmos w=2u l=1u
M6143 n3460 net1854 VSS VSS nmos w=1u l=1u
M6144 net1854 n3462 VSS VSS nmos w=1u l=1u
M6145 net1854 n3463 VSS VSS nmos w=1u l=1u
M6146 net1854 n3463 net1855 VDD pmos w=2u l=1u
M6147 n3460 net1854 VDD VDD pmos w=2u l=1u
M6148 net1855 n3462 VDD VDD pmos w=2u l=1u
M6149 net1856 n3306 VSS VSS nmos w=1u l=1u
M6150 net1857 n3307 VSS VSS nmos w=1u l=1u
M6151 n3458 net1858 VSS VSS nmos w=1u l=1u
M6152 net1858 n3306 net1859 VSS nmos w=1u l=1u
M6153 net1858 net1856 net1857 VSS nmos w=1u l=1u
M6154 net1859 net1857 VSS VSS nmos w=1u l=1u
M6155 net1858 net1856 net1860 VDD pmos w=2u l=1u
M6156 net1856 n3306 VDD VDD pmos w=2u l=1u
M6157 net1857 n3306 net1858 VDD pmos w=2u l=1u
M6158 net1857 n3307 VDD VDD pmos w=2u l=1u
M6159 n3458 net1858 VDD VDD pmos w=2u l=1u
M6160 net1860 net1857 VDD VDD pmos w=2u l=1u
M6161 n3307 n3464 VDD VDD pmos w=2u l=1u
M6162 n3307 n3464 VSS VSS nmos w=1u l=1u
M6163 n3457 n3466 net1861 VSS nmos w=1u l=1u
M6164 net1861 n3465 VSS VSS nmos w=1u l=1u
M6165 n3457 n3466 VDD VDD pmos w=2u l=1u
M6166 n3457 n3465 VDD VDD pmos w=2u l=1u
M6167 net1862 n3464 VSS VSS nmos w=1u l=1u
M6168 net1863 n3306 VSS VSS nmos w=1u l=1u
M6169 n3466 net1864 VSS VSS nmos w=1u l=1u
M6170 net1864 n3464 net1865 VSS nmos w=1u l=1u
M6171 net1864 net1862 net1863 VSS nmos w=1u l=1u
M6172 net1865 net1863 VSS VSS nmos w=1u l=1u
M6173 net1864 net1862 net1866 VDD pmos w=2u l=1u
M6174 net1862 n3464 VDD VDD pmos w=2u l=1u
M6175 net1863 n3464 net1864 VDD pmos w=2u l=1u
M6176 net1863 n3306 VDD VDD pmos w=2u l=1u
M6177 n3466 net1864 VDD VDD pmos w=2u l=1u
M6178 net1866 net1863 VDD VDD pmos w=2u l=1u
M6179 n3464 N494 net1867 VSS nmos w=1u l=1u
M6180 net1867 N52 VSS VSS nmos w=1u l=1u
M6181 n3464 N494 VDD VDD pmos w=2u l=1u
M6182 n3464 N52 VDD VDD pmos w=2u l=1u
M6183 n3306 n3305 net1868 VSS nmos w=1u l=1u
M6184 net1868 n3467 VSS VSS nmos w=1u l=1u
M6185 n3306 n3305 VDD VDD pmos w=2u l=1u
M6186 n3306 n3467 VDD VDD pmos w=2u l=1u
M6187 n3305 n3469 net1869 VSS nmos w=1u l=1u
M6188 net1869 n3468 VSS VSS nmos w=1u l=1u
M6189 n3305 n3469 VDD VDD pmos w=2u l=1u
M6190 n3305 n3468 VDD VDD pmos w=2u l=1u
M6191 n3469 n3471 net1870 VSS nmos w=1u l=1u
M6192 net1870 n3470 VSS VSS nmos w=1u l=1u
M6193 n3469 n3471 VDD VDD pmos w=2u l=1u
M6194 n3469 n3470 VDD VDD pmos w=2u l=1u
M6195 n3470 net1871 VSS VSS nmos w=1u l=1u
M6196 net1871 n3472 VSS VSS nmos w=1u l=1u
M6197 net1871 n3473 VSS VSS nmos w=1u l=1u
M6198 net1871 n3473 net1872 VDD pmos w=2u l=1u
M6199 n3470 net1871 VDD VDD pmos w=2u l=1u
M6200 net1872 n3472 VDD VDD pmos w=2u l=1u
M6201 net1873 n3316 VSS VSS nmos w=1u l=1u
M6202 net1874 n3317 VSS VSS nmos w=1u l=1u
M6203 n3468 net1875 VSS VSS nmos w=1u l=1u
M6204 net1875 n3316 net1876 VSS nmos w=1u l=1u
M6205 net1875 net1873 net1874 VSS nmos w=1u l=1u
M6206 net1876 net1874 VSS VSS nmos w=1u l=1u
M6207 net1875 net1873 net1877 VDD pmos w=2u l=1u
M6208 net1873 n3316 VDD VDD pmos w=2u l=1u
M6209 net1874 n3316 net1875 VDD pmos w=2u l=1u
M6210 net1874 n3317 VDD VDD pmos w=2u l=1u
M6211 n3468 net1875 VDD VDD pmos w=2u l=1u
M6212 net1877 net1874 VDD VDD pmos w=2u l=1u
M6213 n3317 n3474 VDD VDD pmos w=2u l=1u
M6214 n3317 n3474 VSS VSS nmos w=1u l=1u
M6215 n3467 n3476 net1878 VSS nmos w=1u l=1u
M6216 net1878 n3475 VSS VSS nmos w=1u l=1u
M6217 n3467 n3476 VDD VDD pmos w=2u l=1u
M6218 n3467 n3475 VDD VDD pmos w=2u l=1u
M6219 net1879 n3474 VSS VSS nmos w=1u l=1u
M6220 net1880 n3316 VSS VSS nmos w=1u l=1u
M6221 n3476 net1881 VSS VSS nmos w=1u l=1u
M6222 net1881 n3474 net1882 VSS nmos w=1u l=1u
M6223 net1881 net1879 net1880 VSS nmos w=1u l=1u
M6224 net1882 net1880 VSS VSS nmos w=1u l=1u
M6225 net1881 net1879 net1883 VDD pmos w=2u l=1u
M6226 net1879 n3474 VDD VDD pmos w=2u l=1u
M6227 net1880 n3474 net1881 VDD pmos w=2u l=1u
M6228 net1880 n3316 VDD VDD pmos w=2u l=1u
M6229 n3476 net1881 VDD VDD pmos w=2u l=1u
M6230 net1883 net1880 VDD VDD pmos w=2u l=1u
M6231 n3474 N477 net1884 VSS nmos w=1u l=1u
M6232 net1884 N69 VSS VSS nmos w=1u l=1u
M6233 n3474 N477 VDD VDD pmos w=2u l=1u
M6234 n3474 N69 VDD VDD pmos w=2u l=1u
M6235 n3316 n3315 net1885 VSS nmos w=1u l=1u
M6236 net1885 n3477 VSS VSS nmos w=1u l=1u
M6237 n3316 n3315 VDD VDD pmos w=2u l=1u
M6238 n3316 n3477 VDD VDD pmos w=2u l=1u
M6239 n3315 n3479 net1886 VSS nmos w=1u l=1u
M6240 net1886 n3478 VSS VSS nmos w=1u l=1u
M6241 n3315 n3479 VDD VDD pmos w=2u l=1u
M6242 n3315 n3478 VDD VDD pmos w=2u l=1u
M6243 n3479 n3481 net1887 VSS nmos w=1u l=1u
M6244 net1887 n3480 VSS VSS nmos w=1u l=1u
M6245 n3479 n3481 VDD VDD pmos w=2u l=1u
M6246 n3479 n3480 VDD VDD pmos w=2u l=1u
M6247 n3480 net1888 VSS VSS nmos w=1u l=1u
M6248 net1888 n3482 VSS VSS nmos w=1u l=1u
M6249 net1888 n3483 VSS VSS nmos w=1u l=1u
M6250 net1888 n3483 net1889 VDD pmos w=2u l=1u
M6251 n3480 net1888 VDD VDD pmos w=2u l=1u
M6252 net1889 n3482 VDD VDD pmos w=2u l=1u
M6253 net1890 n3326 VSS VSS nmos w=1u l=1u
M6254 net1891 n3327 VSS VSS nmos w=1u l=1u
M6255 n3478 net1892 VSS VSS nmos w=1u l=1u
M6256 net1892 n3326 net1893 VSS nmos w=1u l=1u
M6257 net1892 net1890 net1891 VSS nmos w=1u l=1u
M6258 net1893 net1891 VSS VSS nmos w=1u l=1u
M6259 net1892 net1890 net1894 VDD pmos w=2u l=1u
M6260 net1890 n3326 VDD VDD pmos w=2u l=1u
M6261 net1891 n3326 net1892 VDD pmos w=2u l=1u
M6262 net1891 n3327 VDD VDD pmos w=2u l=1u
M6263 n3478 net1892 VDD VDD pmos w=2u l=1u
M6264 net1894 net1891 VDD VDD pmos w=2u l=1u
M6265 n3327 n3484 VDD VDD pmos w=2u l=1u
M6266 n3327 n3484 VSS VSS nmos w=1u l=1u
M6267 n3477 n3486 net1895 VSS nmos w=1u l=1u
M6268 net1895 n3485 VSS VSS nmos w=1u l=1u
M6269 n3477 n3486 VDD VDD pmos w=2u l=1u
M6270 n3477 n3485 VDD VDD pmos w=2u l=1u
M6271 net1896 n3484 VSS VSS nmos w=1u l=1u
M6272 net1897 n3326 VSS VSS nmos w=1u l=1u
M6273 n3486 net1898 VSS VSS nmos w=1u l=1u
M6274 net1898 n3484 net1899 VSS nmos w=1u l=1u
M6275 net1898 net1896 net1897 VSS nmos w=1u l=1u
M6276 net1899 net1897 VSS VSS nmos w=1u l=1u
M6277 net1898 net1896 net1900 VDD pmos w=2u l=1u
M6278 net1896 n3484 VDD VDD pmos w=2u l=1u
M6279 net1897 n3484 net1898 VDD pmos w=2u l=1u
M6280 net1897 n3326 VDD VDD pmos w=2u l=1u
M6281 n3486 net1898 VDD VDD pmos w=2u l=1u
M6282 net1900 net1897 VDD VDD pmos w=2u l=1u
M6283 n3484 N460 net1901 VSS nmos w=1u l=1u
M6284 net1901 N86 VSS VSS nmos w=1u l=1u
M6285 n3484 N460 VDD VDD pmos w=2u l=1u
M6286 n3484 N86 VDD VDD pmos w=2u l=1u
M6287 n3326 n3325 net1902 VSS nmos w=1u l=1u
M6288 net1902 n3487 VSS VSS nmos w=1u l=1u
M6289 n3326 n3325 VDD VDD pmos w=2u l=1u
M6290 n3326 n3487 VDD VDD pmos w=2u l=1u
M6291 n3325 n3489 net1903 VSS nmos w=1u l=1u
M6292 net1903 n3488 VSS VSS nmos w=1u l=1u
M6293 n3325 n3489 VDD VDD pmos w=2u l=1u
M6294 n3325 n3488 VDD VDD pmos w=2u l=1u
M6295 n3489 n3491 net1904 VSS nmos w=1u l=1u
M6296 net1904 n3490 VSS VSS nmos w=1u l=1u
M6297 n3489 n3491 VDD VDD pmos w=2u l=1u
M6298 n3489 n3490 VDD VDD pmos w=2u l=1u
M6299 n3490 net1905 VSS VSS nmos w=1u l=1u
M6300 net1905 n3492 VSS VSS nmos w=1u l=1u
M6301 net1905 n3493 VSS VSS nmos w=1u l=1u
M6302 net1905 n3493 net1906 VDD pmos w=2u l=1u
M6303 n3490 net1905 VDD VDD pmos w=2u l=1u
M6304 net1906 n3492 VDD VDD pmos w=2u l=1u
M6305 net1907 n3336 VSS VSS nmos w=1u l=1u
M6306 net1908 n3337 VSS VSS nmos w=1u l=1u
M6307 n3488 net1909 VSS VSS nmos w=1u l=1u
M6308 net1909 n3336 net1910 VSS nmos w=1u l=1u
M6309 net1909 net1907 net1908 VSS nmos w=1u l=1u
M6310 net1910 net1908 VSS VSS nmos w=1u l=1u
M6311 net1909 net1907 net1911 VDD pmos w=2u l=1u
M6312 net1907 n3336 VDD VDD pmos w=2u l=1u
M6313 net1908 n3336 net1909 VDD pmos w=2u l=1u
M6314 net1908 n3337 VDD VDD pmos w=2u l=1u
M6315 n3488 net1909 VDD VDD pmos w=2u l=1u
M6316 net1911 net1908 VDD VDD pmos w=2u l=1u
M6317 n3337 n3494 VDD VDD pmos w=2u l=1u
M6318 n3337 n3494 VSS VSS nmos w=1u l=1u
M6319 n3487 n3496 net1912 VSS nmos w=1u l=1u
M6320 net1912 n3495 VSS VSS nmos w=1u l=1u
M6321 n3487 n3496 VDD VDD pmos w=2u l=1u
M6322 n3487 n3495 VDD VDD pmos w=2u l=1u
M6323 net1913 n3494 VSS VSS nmos w=1u l=1u
M6324 net1914 n3336 VSS VSS nmos w=1u l=1u
M6325 n3496 net1915 VSS VSS nmos w=1u l=1u
M6326 net1915 n3494 net1916 VSS nmos w=1u l=1u
M6327 net1915 net1913 net1914 VSS nmos w=1u l=1u
M6328 net1916 net1914 VSS VSS nmos w=1u l=1u
M6329 net1915 net1913 net1917 VDD pmos w=2u l=1u
M6330 net1913 n3494 VDD VDD pmos w=2u l=1u
M6331 net1914 n3494 net1915 VDD pmos w=2u l=1u
M6332 net1914 n3336 VDD VDD pmos w=2u l=1u
M6333 n3496 net1915 VDD VDD pmos w=2u l=1u
M6334 net1917 net1914 VDD VDD pmos w=2u l=1u
M6335 n3494 N443 net1918 VSS nmos w=1u l=1u
M6336 net1918 N103 VSS VSS nmos w=1u l=1u
M6337 n3494 N443 VDD VDD pmos w=2u l=1u
M6338 n3494 N103 VDD VDD pmos w=2u l=1u
M6339 n3336 n3335 net1919 VSS nmos w=1u l=1u
M6340 net1919 n3497 VSS VSS nmos w=1u l=1u
M6341 n3336 n3335 VDD VDD pmos w=2u l=1u
M6342 n3336 n3497 VDD VDD pmos w=2u l=1u
M6343 n3335 n3499 net1920 VSS nmos w=1u l=1u
M6344 net1920 n3498 VSS VSS nmos w=1u l=1u
M6345 n3335 n3499 VDD VDD pmos w=2u l=1u
M6346 n3335 n3498 VDD VDD pmos w=2u l=1u
M6347 n3499 n3501 net1921 VSS nmos w=1u l=1u
M6348 net1921 n3500 VSS VSS nmos w=1u l=1u
M6349 n3499 n3501 VDD VDD pmos w=2u l=1u
M6350 n3499 n3500 VDD VDD pmos w=2u l=1u
M6351 n3500 net1922 VSS VSS nmos w=1u l=1u
M6352 net1922 n3502 VSS VSS nmos w=1u l=1u
M6353 net1922 n3503 VSS VSS nmos w=1u l=1u
M6354 net1922 n3503 net1923 VDD pmos w=2u l=1u
M6355 n3500 net1922 VDD VDD pmos w=2u l=1u
M6356 net1923 n3502 VDD VDD pmos w=2u l=1u
M6357 net1924 n3346 VSS VSS nmos w=1u l=1u
M6358 net1925 n3347 VSS VSS nmos w=1u l=1u
M6359 n3498 net1926 VSS VSS nmos w=1u l=1u
M6360 net1926 n3346 net1927 VSS nmos w=1u l=1u
M6361 net1926 net1924 net1925 VSS nmos w=1u l=1u
M6362 net1927 net1925 VSS VSS nmos w=1u l=1u
M6363 net1926 net1924 net1928 VDD pmos w=2u l=1u
M6364 net1924 n3346 VDD VDD pmos w=2u l=1u
M6365 net1925 n3346 net1926 VDD pmos w=2u l=1u
M6366 net1925 n3347 VDD VDD pmos w=2u l=1u
M6367 n3498 net1926 VDD VDD pmos w=2u l=1u
M6368 net1928 net1925 VDD VDD pmos w=2u l=1u
M6369 n3347 n3504 VDD VDD pmos w=2u l=1u
M6370 n3347 n3504 VSS VSS nmos w=1u l=1u
M6371 n3497 n3506 net1929 VSS nmos w=1u l=1u
M6372 net1929 n3505 VSS VSS nmos w=1u l=1u
M6373 n3497 n3506 VDD VDD pmos w=2u l=1u
M6374 n3497 n3505 VDD VDD pmos w=2u l=1u
M6375 net1930 n3504 VSS VSS nmos w=1u l=1u
M6376 net1931 n3346 VSS VSS nmos w=1u l=1u
M6377 n3506 net1932 VSS VSS nmos w=1u l=1u
M6378 net1932 n3504 net1933 VSS nmos w=1u l=1u
M6379 net1932 net1930 net1931 VSS nmos w=1u l=1u
M6380 net1933 net1931 VSS VSS nmos w=1u l=1u
M6381 net1932 net1930 net1934 VDD pmos w=2u l=1u
M6382 net1930 n3504 VDD VDD pmos w=2u l=1u
M6383 net1931 n3504 net1932 VDD pmos w=2u l=1u
M6384 net1931 n3346 VDD VDD pmos w=2u l=1u
M6385 n3506 net1932 VDD VDD pmos w=2u l=1u
M6386 net1934 net1931 VDD VDD pmos w=2u l=1u
M6387 n3504 N426 net1935 VSS nmos w=1u l=1u
M6388 net1935 N120 VSS VSS nmos w=1u l=1u
M6389 n3504 N426 VDD VDD pmos w=2u l=1u
M6390 n3504 N120 VDD VDD pmos w=2u l=1u
M6391 n3346 n3345 net1936 VSS nmos w=1u l=1u
M6392 net1936 n3507 VSS VSS nmos w=1u l=1u
M6393 n3346 n3345 VDD VDD pmos w=2u l=1u
M6394 n3346 n3507 VDD VDD pmos w=2u l=1u
M6395 n3345 n3509 net1937 VSS nmos w=1u l=1u
M6396 net1937 n3508 VSS VSS nmos w=1u l=1u
M6397 n3345 n3509 VDD VDD pmos w=2u l=1u
M6398 n3345 n3508 VDD VDD pmos w=2u l=1u
M6399 n3509 n3511 net1938 VSS nmos w=1u l=1u
M6400 net1938 n3510 VSS VSS nmos w=1u l=1u
M6401 n3509 n3511 VDD VDD pmos w=2u l=1u
M6402 n3509 n3510 VDD VDD pmos w=2u l=1u
M6403 n3510 net1939 VSS VSS nmos w=1u l=1u
M6404 net1939 n3512 VSS VSS nmos w=1u l=1u
M6405 net1939 n3513 VSS VSS nmos w=1u l=1u
M6406 net1939 n3513 net1940 VDD pmos w=2u l=1u
M6407 n3510 net1939 VDD VDD pmos w=2u l=1u
M6408 net1940 n3512 VDD VDD pmos w=2u l=1u
M6409 net1941 n3356 VSS VSS nmos w=1u l=1u
M6410 net1942 n3357 VSS VSS nmos w=1u l=1u
M6411 n3508 net1943 VSS VSS nmos w=1u l=1u
M6412 net1943 n3356 net1944 VSS nmos w=1u l=1u
M6413 net1943 net1941 net1942 VSS nmos w=1u l=1u
M6414 net1944 net1942 VSS VSS nmos w=1u l=1u
M6415 net1943 net1941 net1945 VDD pmos w=2u l=1u
M6416 net1941 n3356 VDD VDD pmos w=2u l=1u
M6417 net1942 n3356 net1943 VDD pmos w=2u l=1u
M6418 net1942 n3357 VDD VDD pmos w=2u l=1u
M6419 n3508 net1943 VDD VDD pmos w=2u l=1u
M6420 net1945 net1942 VDD VDD pmos w=2u l=1u
M6421 n3357 n3514 VDD VDD pmos w=2u l=1u
M6422 n3357 n3514 VSS VSS nmos w=1u l=1u
M6423 n3507 n3516 net1946 VSS nmos w=1u l=1u
M6424 net1946 n3515 VSS VSS nmos w=1u l=1u
M6425 n3507 n3516 VDD VDD pmos w=2u l=1u
M6426 n3507 n3515 VDD VDD pmos w=2u l=1u
M6427 net1947 n3514 VSS VSS nmos w=1u l=1u
M6428 net1948 n3356 VSS VSS nmos w=1u l=1u
M6429 n3516 net1949 VSS VSS nmos w=1u l=1u
M6430 net1949 n3514 net1950 VSS nmos w=1u l=1u
M6431 net1949 net1947 net1948 VSS nmos w=1u l=1u
M6432 net1950 net1948 VSS VSS nmos w=1u l=1u
M6433 net1949 net1947 net1951 VDD pmos w=2u l=1u
M6434 net1947 n3514 VDD VDD pmos w=2u l=1u
M6435 net1948 n3514 net1949 VDD pmos w=2u l=1u
M6436 net1948 n3356 VDD VDD pmos w=2u l=1u
M6437 n3516 net1949 VDD VDD pmos w=2u l=1u
M6438 net1951 net1948 VDD VDD pmos w=2u l=1u
M6439 n3514 N409 net1952 VSS nmos w=1u l=1u
M6440 net1952 N137 VSS VSS nmos w=1u l=1u
M6441 n3514 N409 VDD VDD pmos w=2u l=1u
M6442 n3514 N137 VDD VDD pmos w=2u l=1u
M6443 n3356 n3355 net1953 VSS nmos w=1u l=1u
M6444 net1953 n3517 VSS VSS nmos w=1u l=1u
M6445 n3356 n3355 VDD VDD pmos w=2u l=1u
M6446 n3356 n3517 VDD VDD pmos w=2u l=1u
M6447 n3355 n3519 net1954 VSS nmos w=1u l=1u
M6448 net1954 n3518 VSS VSS nmos w=1u l=1u
M6449 n3355 n3519 VDD VDD pmos w=2u l=1u
M6450 n3355 n3518 VDD VDD pmos w=2u l=1u
M6451 n3519 n3521 net1955 VSS nmos w=1u l=1u
M6452 net1955 n3520 VSS VSS nmos w=1u l=1u
M6453 n3519 n3521 VDD VDD pmos w=2u l=1u
M6454 n3519 n3520 VDD VDD pmos w=2u l=1u
M6455 n3520 net1956 VSS VSS nmos w=1u l=1u
M6456 net1956 n3522 VSS VSS nmos w=1u l=1u
M6457 net1956 n3523 VSS VSS nmos w=1u l=1u
M6458 net1956 n3523 net1957 VDD pmos w=2u l=1u
M6459 n3520 net1956 VDD VDD pmos w=2u l=1u
M6460 net1957 n3522 VDD VDD pmos w=2u l=1u
M6461 net1958 n3366 VSS VSS nmos w=1u l=1u
M6462 net1959 n3367 VSS VSS nmos w=1u l=1u
M6463 n3518 net1960 VSS VSS nmos w=1u l=1u
M6464 net1960 n3366 net1961 VSS nmos w=1u l=1u
M6465 net1960 net1958 net1959 VSS nmos w=1u l=1u
M6466 net1961 net1959 VSS VSS nmos w=1u l=1u
M6467 net1960 net1958 net1962 VDD pmos w=2u l=1u
M6468 net1958 n3366 VDD VDD pmos w=2u l=1u
M6469 net1959 n3366 net1960 VDD pmos w=2u l=1u
M6470 net1959 n3367 VDD VDD pmos w=2u l=1u
M6471 n3518 net1960 VDD VDD pmos w=2u l=1u
M6472 net1962 net1959 VDD VDD pmos w=2u l=1u
M6473 n3367 n3524 VDD VDD pmos w=2u l=1u
M6474 n3367 n3524 VSS VSS nmos w=1u l=1u
M6475 n3517 n3526 net1963 VSS nmos w=1u l=1u
M6476 net1963 n3525 VSS VSS nmos w=1u l=1u
M6477 n3517 n3526 VDD VDD pmos w=2u l=1u
M6478 n3517 n3525 VDD VDD pmos w=2u l=1u
M6479 net1964 n3524 VSS VSS nmos w=1u l=1u
M6480 net1965 n3366 VSS VSS nmos w=1u l=1u
M6481 n3526 net1966 VSS VSS nmos w=1u l=1u
M6482 net1966 n3524 net1967 VSS nmos w=1u l=1u
M6483 net1966 net1964 net1965 VSS nmos w=1u l=1u
M6484 net1967 net1965 VSS VSS nmos w=1u l=1u
M6485 net1966 net1964 net1968 VDD pmos w=2u l=1u
M6486 net1964 n3524 VDD VDD pmos w=2u l=1u
M6487 net1965 n3524 net1966 VDD pmos w=2u l=1u
M6488 net1965 n3366 VDD VDD pmos w=2u l=1u
M6489 n3526 net1966 VDD VDD pmos w=2u l=1u
M6490 net1968 net1965 VDD VDD pmos w=2u l=1u
M6491 n3524 N392 net1969 VSS nmos w=1u l=1u
M6492 net1969 N154 VSS VSS nmos w=1u l=1u
M6493 n3524 N392 VDD VDD pmos w=2u l=1u
M6494 n3524 N154 VDD VDD pmos w=2u l=1u
M6495 n3366 n3365 net1970 VSS nmos w=1u l=1u
M6496 net1970 n3527 VSS VSS nmos w=1u l=1u
M6497 n3366 n3365 VDD VDD pmos w=2u l=1u
M6498 n3366 n3527 VDD VDD pmos w=2u l=1u
M6499 n3365 n3529 net1971 VSS nmos w=1u l=1u
M6500 net1971 n3528 VSS VSS nmos w=1u l=1u
M6501 n3365 n3529 VDD VDD pmos w=2u l=1u
M6502 n3365 n3528 VDD VDD pmos w=2u l=1u
M6503 n3529 n3531 net1972 VSS nmos w=1u l=1u
M6504 net1972 n3530 VSS VSS nmos w=1u l=1u
M6505 n3529 n3531 VDD VDD pmos w=2u l=1u
M6506 n3529 n3530 VDD VDD pmos w=2u l=1u
M6507 n3530 n3533 net1973 VSS nmos w=1u l=1u
M6508 net1973 n3532 VSS VSS nmos w=1u l=1u
M6509 n3530 n3533 VDD VDD pmos w=2u l=1u
M6510 n3530 n3532 VDD VDD pmos w=2u l=1u
M6511 net1974 n3376 VSS VSS nmos w=1u l=1u
M6512 net1975 n3377 VSS VSS nmos w=1u l=1u
M6513 n3528 net1976 VSS VSS nmos w=1u l=1u
M6514 net1976 n3376 net1977 VSS nmos w=1u l=1u
M6515 net1976 net1974 net1975 VSS nmos w=1u l=1u
M6516 net1977 net1975 VSS VSS nmos w=1u l=1u
M6517 net1976 net1974 net1978 VDD pmos w=2u l=1u
M6518 net1974 n3376 VDD VDD pmos w=2u l=1u
M6519 net1975 n3376 net1976 VDD pmos w=2u l=1u
M6520 net1975 n3377 VDD VDD pmos w=2u l=1u
M6521 n3528 net1976 VDD VDD pmos w=2u l=1u
M6522 net1978 net1975 VDD VDD pmos w=2u l=1u
M6523 n3376 n3534 VDD VDD pmos w=2u l=1u
M6524 n3376 n3534 VSS VSS nmos w=1u l=1u
M6525 n3527 n3536 net1979 VSS nmos w=1u l=1u
M6526 net1979 n3535 VSS VSS nmos w=1u l=1u
M6527 n3527 n3536 VDD VDD pmos w=2u l=1u
M6528 n3527 n3535 VDD VDD pmos w=2u l=1u
M6529 net1980 n3377 VSS VSS nmos w=1u l=1u
M6530 net1981 n3534 VSS VSS nmos w=1u l=1u
M6531 n3536 net1982 VSS VSS nmos w=1u l=1u
M6532 net1982 n3377 net1983 VSS nmos w=1u l=1u
M6533 net1982 net1980 net1981 VSS nmos w=1u l=1u
M6534 net1983 net1981 VSS VSS nmos w=1u l=1u
M6535 net1982 net1980 net1984 VDD pmos w=2u l=1u
M6536 net1980 n3377 VDD VDD pmos w=2u l=1u
M6537 net1981 n3377 net1982 VDD pmos w=2u l=1u
M6538 net1981 n3534 VDD VDD pmos w=2u l=1u
M6539 n3536 net1982 VDD VDD pmos w=2u l=1u
M6540 net1984 net1981 VDD VDD pmos w=2u l=1u
M6541 n3377 N375 net1985 VSS nmos w=1u l=1u
M6542 net1985 N171 VSS VSS nmos w=1u l=1u
M6543 n3377 N375 VDD VDD pmos w=2u l=1u
M6544 n3377 N171 VDD VDD pmos w=2u l=1u
M6545 n3534 n3375 net1986 VSS nmos w=1u l=1u
M6546 net1986 n3537 VSS VSS nmos w=1u l=1u
M6547 n3534 n3375 VDD VDD pmos w=2u l=1u
M6548 n3534 n3537 VDD VDD pmos w=2u l=1u
M6549 n3375 n3539 net1987 VSS nmos w=1u l=1u
M6550 net1987 n3538 VSS VSS nmos w=1u l=1u
M6551 n3375 n3539 VDD VDD pmos w=2u l=1u
M6552 n3375 n3538 VDD VDD pmos w=2u l=1u
M6553 n3539 n3541 net1988 VSS nmos w=1u l=1u
M6554 net1988 n3540 VSS VSS nmos w=1u l=1u
M6555 n3539 n3541 VDD VDD pmos w=2u l=1u
M6556 n3539 n3540 VDD VDD pmos w=2u l=1u
M6557 n3540 net1989 VSS VSS nmos w=1u l=1u
M6558 net1989 n3542 VSS VSS nmos w=1u l=1u
M6559 net1989 n3543 VSS VSS nmos w=1u l=1u
M6560 net1989 n3543 net1990 VDD pmos w=2u l=1u
M6561 n3540 net1989 VDD VDD pmos w=2u l=1u
M6562 net1990 n3542 VDD VDD pmos w=2u l=1u
M6563 net1991 n3386 VSS VSS nmos w=1u l=1u
M6564 net1992 n3387 VSS VSS nmos w=1u l=1u
M6565 n3538 net1993 VSS VSS nmos w=1u l=1u
M6566 net1993 n3386 net1994 VSS nmos w=1u l=1u
M6567 net1993 net1991 net1992 VSS nmos w=1u l=1u
M6568 net1994 net1992 VSS VSS nmos w=1u l=1u
M6569 net1993 net1991 net1995 VDD pmos w=2u l=1u
M6570 net1991 n3386 VDD VDD pmos w=2u l=1u
M6571 net1992 n3386 net1993 VDD pmos w=2u l=1u
M6572 net1992 n3387 VDD VDD pmos w=2u l=1u
M6573 n3538 net1993 VDD VDD pmos w=2u l=1u
M6574 net1995 net1992 VDD VDD pmos w=2u l=1u
M6575 n3387 n3544 VDD VDD pmos w=2u l=1u
M6576 n3387 n3544 VSS VSS nmos w=1u l=1u
M6577 n3537 n3546 net1996 VSS nmos w=1u l=1u
M6578 net1996 n3545 VSS VSS nmos w=1u l=1u
M6579 n3537 n3546 VDD VDD pmos w=2u l=1u
M6580 n3537 n3545 VDD VDD pmos w=2u l=1u
M6581 net1997 n3544 VSS VSS nmos w=1u l=1u
M6582 net1998 n3386 VSS VSS nmos w=1u l=1u
M6583 n3546 net1999 VSS VSS nmos w=1u l=1u
M6584 net1999 n3544 net2000 VSS nmos w=1u l=1u
M6585 net1999 net1997 net1998 VSS nmos w=1u l=1u
M6586 net2000 net1998 VSS VSS nmos w=1u l=1u
M6587 net1999 net1997 net2001 VDD pmos w=2u l=1u
M6588 net1997 n3544 VDD VDD pmos w=2u l=1u
M6589 net1998 n3544 net1999 VDD pmos w=2u l=1u
M6590 net1998 n3386 VDD VDD pmos w=2u l=1u
M6591 n3546 net1999 VDD VDD pmos w=2u l=1u
M6592 net2001 net1998 VDD VDD pmos w=2u l=1u
M6593 n3544 N358 net2002 VSS nmos w=1u l=1u
M6594 net2002 N188 VSS VSS nmos w=1u l=1u
M6595 n3544 N358 VDD VDD pmos w=2u l=1u
M6596 n3544 N188 VDD VDD pmos w=2u l=1u
M6597 n3386 n3385 net2003 VSS nmos w=1u l=1u
M6598 net2003 n3547 VSS VSS nmos w=1u l=1u
M6599 n3386 n3385 VDD VDD pmos w=2u l=1u
M6600 n3386 n3547 VDD VDD pmos w=2u l=1u
M6601 n3385 n3549 net2004 VSS nmos w=1u l=1u
M6602 net2004 n3548 VSS VSS nmos w=1u l=1u
M6603 n3385 n3549 VDD VDD pmos w=2u l=1u
M6604 n3385 n3548 VDD VDD pmos w=2u l=1u
M6605 n3549 n3551 net2005 VSS nmos w=1u l=1u
M6606 net2005 n3550 VSS VSS nmos w=1u l=1u
M6607 n3549 n3551 VDD VDD pmos w=2u l=1u
M6608 n3549 n3550 VDD VDD pmos w=2u l=1u
M6609 n3550 net2006 VSS VSS nmos w=1u l=1u
M6610 net2006 n3552 VSS VSS nmos w=1u l=1u
M6611 net2006 n3553 VSS VSS nmos w=1u l=1u
M6612 net2006 n3553 net2007 VDD pmos w=2u l=1u
M6613 n3550 net2006 VDD VDD pmos w=2u l=1u
M6614 net2007 n3552 VDD VDD pmos w=2u l=1u
M6615 net2008 n3396 VSS VSS nmos w=1u l=1u
M6616 net2009 n3397 VSS VSS nmos w=1u l=1u
M6617 n3548 net2010 VSS VSS nmos w=1u l=1u
M6618 net2010 n3396 net2011 VSS nmos w=1u l=1u
M6619 net2010 net2008 net2009 VSS nmos w=1u l=1u
M6620 net2011 net2009 VSS VSS nmos w=1u l=1u
M6621 net2010 net2008 net2012 VDD pmos w=2u l=1u
M6622 net2008 n3396 VDD VDD pmos w=2u l=1u
M6623 net2009 n3396 net2010 VDD pmos w=2u l=1u
M6624 net2009 n3397 VDD VDD pmos w=2u l=1u
M6625 n3548 net2010 VDD VDD pmos w=2u l=1u
M6626 net2012 net2009 VDD VDD pmos w=2u l=1u
M6627 n3397 n3554 VDD VDD pmos w=2u l=1u
M6628 n3397 n3554 VSS VSS nmos w=1u l=1u
M6629 n3547 n3556 net2013 VSS nmos w=1u l=1u
M6630 net2013 n3555 VSS VSS nmos w=1u l=1u
M6631 n3547 n3556 VDD VDD pmos w=2u l=1u
M6632 n3547 n3555 VDD VDD pmos w=2u l=1u
M6633 net2014 n3554 VSS VSS nmos w=1u l=1u
M6634 net2015 n3396 VSS VSS nmos w=1u l=1u
M6635 n3556 net2016 VSS VSS nmos w=1u l=1u
M6636 net2016 n3554 net2017 VSS nmos w=1u l=1u
M6637 net2016 net2014 net2015 VSS nmos w=1u l=1u
M6638 net2017 net2015 VSS VSS nmos w=1u l=1u
M6639 net2016 net2014 net2018 VDD pmos w=2u l=1u
M6640 net2014 n3554 VDD VDD pmos w=2u l=1u
M6641 net2015 n3554 net2016 VDD pmos w=2u l=1u
M6642 net2015 n3396 VDD VDD pmos w=2u l=1u
M6643 n3556 net2016 VDD VDD pmos w=2u l=1u
M6644 net2018 net2015 VDD VDD pmos w=2u l=1u
M6645 n3554 N341 net2019 VSS nmos w=1u l=1u
M6646 net2019 N205 VSS VSS nmos w=1u l=1u
M6647 n3554 N341 VDD VDD pmos w=2u l=1u
M6648 n3554 N205 VDD VDD pmos w=2u l=1u
M6649 n3396 n3395 net2020 VSS nmos w=1u l=1u
M6650 net2020 n3557 VSS VSS nmos w=1u l=1u
M6651 n3396 n3395 VDD VDD pmos w=2u l=1u
M6652 n3396 n3557 VDD VDD pmos w=2u l=1u
M6653 n3395 n3559 net2021 VSS nmos w=1u l=1u
M6654 net2021 n3558 VSS VSS nmos w=1u l=1u
M6655 n3395 n3559 VDD VDD pmos w=2u l=1u
M6656 n3395 n3558 VDD VDD pmos w=2u l=1u
M6657 n3559 net2022 VSS VSS nmos w=1u l=1u
M6658 net2022 n3560 VSS VSS nmos w=1u l=1u
M6659 net2022 n3561 VSS VSS nmos w=1u l=1u
M6660 net2022 n3561 net2023 VDD pmos w=2u l=1u
M6661 n3559 net2022 VDD VDD pmos w=2u l=1u
M6662 net2023 n3560 VDD VDD pmos w=2u l=1u
M6663 n3558 net2024 VSS VSS nmos w=1u l=1u
M6664 net2025 n3562 VSS VSS nmos w=1u l=1u
M6665 net2024 n3418 net2025 VSS nmos w=1u l=1u
M6666 net2024 n3562 VDD VDD pmos w=2u l=1u
M6667 net2024 n3418 VDD VDD pmos w=2u l=1u
M6668 n3558 net2024 VDD VDD pmos w=2u l=1u
M6669 n3557 n3564 net2026 VSS nmos w=1u l=1u
M6670 net2026 n3563 VSS VSS nmos w=1u l=1u
M6671 n3557 n3564 VDD VDD pmos w=2u l=1u
M6672 n3557 n3563 VDD VDD pmos w=2u l=1u
M6673 n3564 n3418 net2027 VSS nmos w=1u l=1u
M6674 net2027 n3562 VSS VSS nmos w=1u l=1u
M6675 n3564 n3418 VDD VDD pmos w=2u l=1u
M6676 n3564 n3562 VDD VDD pmos w=2u l=1u
M6677 n3418 n3566 net2028 VSS nmos w=1u l=1u
M6678 net2028 n3565 VSS VSS nmos w=1u l=1u
M6679 n3418 n3566 VDD VDD pmos w=2u l=1u
M6680 n3418 n3565 VDD VDD pmos w=2u l=1u
M6681 n3566 N324 net2029 VSS nmos w=1u l=1u
M6682 net2029 N222 VSS VSS nmos w=1u l=1u
M6683 n3566 N324 VDD VDD pmos w=2u l=1u
M6684 n3566 N222 VDD VDD pmos w=2u l=1u
M6685 n3562 N222 net2030 VSS nmos w=1u l=1u
M6686 net2030 n3567 VSS VSS nmos w=1u l=1u
M6687 n3562 N222 VDD VDD pmos w=2u l=1u
M6688 n3562 n3567 VDD VDD pmos w=2u l=1u
M6689 n3567 n3257 VSS VSS nmos w=1u l=1u
M6690 n3567 n3565 VSS VSS nmos w=1u l=1u
M6691 n3567 n3257 net2031 VDD pmos w=2u l=1u
M6692 net2031 n3565 VDD VDD pmos w=2u l=1u
M6693 n3565 n3416 VSS VSS nmos w=1u l=1u
M6694 n3565 n3568 VSS VSS nmos w=1u l=1u
M6695 n3565 n3416 net2032 VDD pmos w=2u l=1u
M6696 net2032 n3568 VDD VDD pmos w=2u l=1u
M6697 n3416 n3570 VSS VSS nmos w=1u l=1u
M6698 n3416 n3569 VSS VSS nmos w=1u l=1u
M6699 n3416 n3570 net2033 VDD pmos w=2u l=1u
M6700 net2033 n3569 VDD VDD pmos w=2u l=1u
M6701 n3568 net2034 VSS VSS nmos w=1u l=1u
M6702 net2035 n3569 VSS VSS nmos w=1u l=1u
M6703 net2034 n3570 net2035 VSS nmos w=1u l=1u
M6704 net2034 n3569 VDD VDD pmos w=2u l=1u
M6705 net2034 n3570 VDD VDD pmos w=2u l=1u
M6706 n3568 net2034 VDD VDD pmos w=2u l=1u
M6707 n3569 n3571 net2036 VSS nmos w=1u l=1u
M6708 net2036 n3415 VSS VSS nmos w=1u l=1u
M6709 n3569 n3571 VDD VDD pmos w=2u l=1u
M6710 n3569 n3415 VDD VDD pmos w=2u l=1u
M6711 n3571 n3572 net2037 VSS nmos w=1u l=1u
M6712 net2037 N307 VSS VSS nmos w=1u l=1u
M6713 n3571 n3572 VDD VDD pmos w=2u l=1u
M6714 n3571 N307 VDD VDD pmos w=2u l=1u
M6715 n3572 n3573 net2038 VSS nmos w=1u l=1u
M6716 net2038 n2270 VSS VSS nmos w=1u l=1u
M6717 n3572 n3573 VDD VDD pmos w=2u l=1u
M6718 n3572 n2270 VDD VDD pmos w=2u l=1u
M6719 n3573 n3574 net2039 VSS nmos w=1u l=1u
M6720 net2039 N239 VSS VSS nmos w=1u l=1u
M6721 n3573 n3574 VDD VDD pmos w=2u l=1u
M6722 n3573 N239 VDD VDD pmos w=2u l=1u
M6723 n2270 n2275 net2040 VSS nmos w=1u l=1u
M6724 net2040 N239 VSS VSS nmos w=1u l=1u
M6725 n2270 n2275 VDD VDD pmos w=2u l=1u
M6726 n2270 N239 VDD VDD pmos w=2u l=1u
M6727 n3415 n3576 net2041 VSS nmos w=1u l=1u
M6728 net2041 n3575 VSS VSS nmos w=1u l=1u
M6729 n3415 n3576 VDD VDD pmos w=2u l=1u
M6730 n3415 n3575 VDD VDD pmos w=2u l=1u
M6731 n3575 n2275 VSS VSS nmos w=1u l=1u
M6732 n3575 n3577 VSS VSS nmos w=1u l=1u
M6733 n3575 n2275 net2042 VDD pmos w=2u l=1u
M6734 net2042 n3577 VDD VDD pmos w=2u l=1u
M6735 n3577 n3411 VSS VSS nmos w=1u l=1u
M6736 n3577 n2228 VSS VSS nmos w=1u l=1u
M6737 n3577 n3411 net2043 VDD pmos w=2u l=1u
M6738 net2043 n2228 VDD VDD pmos w=2u l=1u
M6739 n3570 net2044 VSS VSS nmos w=1u l=1u
M6740 net2045 n3579 VSS VSS nmos w=1u l=1u
M6741 net2044 n3578 net2045 VSS nmos w=1u l=1u
M6742 net2044 n3579 VDD VDD pmos w=2u l=1u
M6743 net2044 n3578 VDD VDD pmos w=2u l=1u
M6744 n3570 net2044 VDD VDD pmos w=2u l=1u
M6745 n3563 n3560 VSS VSS nmos w=1u l=1u
M6746 n3563 n3561 VSS VSS nmos w=1u l=1u
M6747 n3563 n3560 net2046 VDD pmos w=2u l=1u
M6748 net2046 n3561 VDD VDD pmos w=2u l=1u
M6749 n3560 n3580 VDD VDD pmos w=2u l=1u
M6750 n3560 n3580 VSS VSS nmos w=1u l=1u
M6751 n3555 n3582 VSS VSS nmos w=1u l=1u
M6752 n3555 n3581 VSS VSS nmos w=1u l=1u
M6753 n3555 n3582 net2047 VDD pmos w=2u l=1u
M6754 net2047 n3581 VDD VDD pmos w=2u l=1u
M6755 n3582 n3552 VSS VSS nmos w=1u l=1u
M6756 n3582 n3553 VSS VSS nmos w=1u l=1u
M6757 n3582 n3552 net2048 VDD pmos w=2u l=1u
M6758 net2048 n3553 VDD VDD pmos w=2u l=1u
M6759 n3581 n3551 VDD VDD pmos w=2u l=1u
M6760 n3581 n3551 VSS VSS nmos w=1u l=1u
M6761 n3545 n3584 VSS VSS nmos w=1u l=1u
M6762 n3545 n3583 VSS VSS nmos w=1u l=1u
M6763 n3545 n3584 net2049 VDD pmos w=2u l=1u
M6764 net2049 n3583 VDD VDD pmos w=2u l=1u
M6765 n3584 n3542 VSS VSS nmos w=1u l=1u
M6766 n3584 n3543 VSS VSS nmos w=1u l=1u
M6767 n3584 n3542 net2050 VDD pmos w=2u l=1u
M6768 net2050 n3543 VDD VDD pmos w=2u l=1u
M6769 n3583 n3541 VDD VDD pmos w=2u l=1u
M6770 n3583 n3541 VSS VSS nmos w=1u l=1u
M6771 n3535 n3586 VSS VSS nmos w=1u l=1u
M6772 n3535 n3585 VSS VSS nmos w=1u l=1u
M6773 n3535 n3586 net2051 VDD pmos w=2u l=1u
M6774 net2051 n3585 VDD VDD pmos w=2u l=1u
M6775 n3586 net2052 VSS VSS nmos w=1u l=1u
M6776 net2053 n3532 VSS VSS nmos w=1u l=1u
M6777 net2052 n3533 net2053 VSS nmos w=1u l=1u
M6778 net2052 n3532 VDD VDD pmos w=2u l=1u
M6779 net2052 n3533 VDD VDD pmos w=2u l=1u
M6780 n3586 net2052 VDD VDD pmos w=2u l=1u
M6781 n3585 n3531 VDD VDD pmos w=2u l=1u
M6782 n3585 n3531 VSS VSS nmos w=1u l=1u
M6783 n3525 n3588 VSS VSS nmos w=1u l=1u
M6784 n3525 n3587 VSS VSS nmos w=1u l=1u
M6785 n3525 n3588 net2054 VDD pmos w=2u l=1u
M6786 net2054 n3587 VDD VDD pmos w=2u l=1u
M6787 n3588 n3522 VSS VSS nmos w=1u l=1u
M6788 n3588 n3523 VSS VSS nmos w=1u l=1u
M6789 n3588 n3522 net2055 VDD pmos w=2u l=1u
M6790 net2055 n3523 VDD VDD pmos w=2u l=1u
M6791 n3587 n3521 VDD VDD pmos w=2u l=1u
M6792 n3587 n3521 VSS VSS nmos w=1u l=1u
M6793 n3515 n3590 VSS VSS nmos w=1u l=1u
M6794 n3515 n3589 VSS VSS nmos w=1u l=1u
M6795 n3515 n3590 net2056 VDD pmos w=2u l=1u
M6796 net2056 n3589 VDD VDD pmos w=2u l=1u
M6797 n3590 n3512 VSS VSS nmos w=1u l=1u
M6798 n3590 n3513 VSS VSS nmos w=1u l=1u
M6799 n3590 n3512 net2057 VDD pmos w=2u l=1u
M6800 net2057 n3513 VDD VDD pmos w=2u l=1u
M6801 n3589 n3511 VDD VDD pmos w=2u l=1u
M6802 n3589 n3511 VSS VSS nmos w=1u l=1u
M6803 n3505 n3592 VSS VSS nmos w=1u l=1u
M6804 n3505 n3591 VSS VSS nmos w=1u l=1u
M6805 n3505 n3592 net2058 VDD pmos w=2u l=1u
M6806 net2058 n3591 VDD VDD pmos w=2u l=1u
M6807 n3592 n3502 VSS VSS nmos w=1u l=1u
M6808 n3592 n3503 VSS VSS nmos w=1u l=1u
M6809 n3592 n3502 net2059 VDD pmos w=2u l=1u
M6810 net2059 n3503 VDD VDD pmos w=2u l=1u
M6811 n3591 n3501 VDD VDD pmos w=2u l=1u
M6812 n3591 n3501 VSS VSS nmos w=1u l=1u
M6813 n3495 n3594 VSS VSS nmos w=1u l=1u
M6814 n3495 n3593 VSS VSS nmos w=1u l=1u
M6815 n3495 n3594 net2060 VDD pmos w=2u l=1u
M6816 net2060 n3593 VDD VDD pmos w=2u l=1u
M6817 n3594 n3492 VSS VSS nmos w=1u l=1u
M6818 n3594 n3493 VSS VSS nmos w=1u l=1u
M6819 n3594 n3492 net2061 VDD pmos w=2u l=1u
M6820 net2061 n3493 VDD VDD pmos w=2u l=1u
M6821 n3593 n3491 VDD VDD pmos w=2u l=1u
M6822 n3593 n3491 VSS VSS nmos w=1u l=1u
M6823 n3485 n3596 VSS VSS nmos w=1u l=1u
M6824 n3485 n3595 VSS VSS nmos w=1u l=1u
M6825 n3485 n3596 net2062 VDD pmos w=2u l=1u
M6826 net2062 n3595 VDD VDD pmos w=2u l=1u
M6827 n3596 n3482 VSS VSS nmos w=1u l=1u
M6828 n3596 n3483 VSS VSS nmos w=1u l=1u
M6829 n3596 n3482 net2063 VDD pmos w=2u l=1u
M6830 net2063 n3483 VDD VDD pmos w=2u l=1u
M6831 n3595 n3481 VDD VDD pmos w=2u l=1u
M6832 n3595 n3481 VSS VSS nmos w=1u l=1u
M6833 n3475 n3598 VSS VSS nmos w=1u l=1u
M6834 n3475 n3597 VSS VSS nmos w=1u l=1u
M6835 n3475 n3598 net2064 VDD pmos w=2u l=1u
M6836 net2064 n3597 VDD VDD pmos w=2u l=1u
M6837 n3598 n3472 VSS VSS nmos w=1u l=1u
M6838 n3598 n3473 VSS VSS nmos w=1u l=1u
M6839 n3598 n3472 net2065 VDD pmos w=2u l=1u
M6840 net2065 n3473 VDD VDD pmos w=2u l=1u
M6841 n3597 n3471 VDD VDD pmos w=2u l=1u
M6842 n3597 n3471 VSS VSS nmos w=1u l=1u
M6843 n3465 n3600 VSS VSS nmos w=1u l=1u
M6844 n3465 n3599 VSS VSS nmos w=1u l=1u
M6845 n3465 n3600 net2066 VDD pmos w=2u l=1u
M6846 net2066 n3599 VDD VDD pmos w=2u l=1u
M6847 n3600 n3462 VSS VSS nmos w=1u l=1u
M6848 n3600 n3463 VSS VSS nmos w=1u l=1u
M6849 n3600 n3462 net2067 VDD pmos w=2u l=1u
M6850 net2067 n3463 VDD VDD pmos w=2u l=1u
M6851 n3599 n3461 VDD VDD pmos w=2u l=1u
M6852 n3599 n3461 VSS VSS nmos w=1u l=1u
M6853 n3453 n3602 VSS VSS nmos w=1u l=1u
M6854 n3453 n3601 VSS VSS nmos w=1u l=1u
M6855 n3453 n3602 net2068 VDD pmos w=2u l=1u
M6856 net2068 n3601 VDD VDD pmos w=2u l=1u
M6857 n3602 n3451 VSS VSS nmos w=1u l=1u
M6858 n3602 n3452 VSS VSS nmos w=1u l=1u
M6859 n3602 n3451 net2069 VDD pmos w=2u l=1u
M6860 net2069 n3452 VDD VDD pmos w=2u l=1u
M6861 n3601 n3450 VDD VDD pmos w=2u l=1u
M6862 n3601 n3450 VSS VSS nmos w=1u l=1u
M6863 n3445 n2205 VSS VSS nmos w=1u l=1u
M6864 n3445 n3603 VSS VSS nmos w=1u l=1u
M6865 n3445 n2205 net2070 VDD pmos w=2u l=1u
M6866 net2070 n3603 VDD VDD pmos w=2u l=1u
M6867 n2205 N528 VDD VDD pmos w=2u l=1u
M6868 n2205 N528 VSS VSS nmos w=1u l=1u
M6869 n3443 net2071 VSS VSS nmos w=1u l=1u
M6870 net2072 n3605 VSS VSS nmos w=1u l=1u
M6871 net2071 n3604 net2072 VSS nmos w=1u l=1u
M6872 net2071 n3605 VDD VDD pmos w=2u l=1u
M6873 net2071 n3604 VDD VDD pmos w=2u l=1u
M6874 n3443 net2071 VDD VDD pmos w=2u l=1u
M6875 n3604 n3607 net2073 VSS nmos w=1u l=1u
M6876 net2073 n3606 VSS VSS nmos w=1u l=1u
M6877 n3604 n3607 VDD VDD pmos w=2u l=1u
M6878 n3604 n3606 VDD VDD pmos w=2u l=1u
M6879 n3606 n3608 VDD VDD pmos w=2u l=1u
M6880 n3606 n3608 VSS VSS nmos w=1u l=1u
M6881 net2074 n3607 VSS VSS nmos w=1u l=1u
M6882 net2075 n3608 VSS VSS nmos w=1u l=1u
M6883 N6123 net2076 VSS VSS nmos w=1u l=1u
M6884 net2076 n3607 net2077 VSS nmos w=1u l=1u
M6885 net2076 net2074 net2075 VSS nmos w=1u l=1u
M6886 net2077 net2075 VSS VSS nmos w=1u l=1u
M6887 net2076 net2074 net2078 VDD pmos w=2u l=1u
M6888 net2074 n3607 VDD VDD pmos w=2u l=1u
M6889 net2075 n3607 net2076 VDD pmos w=2u l=1u
M6890 net2075 n3608 VDD VDD pmos w=2u l=1u
M6891 N6123 net2076 VDD VDD pmos w=2u l=1u
M6892 net2078 net2075 VDD VDD pmos w=2u l=1u
M6893 n3607 N528 net2079 VSS nmos w=1u l=1u
M6894 net2079 N1 VSS VSS nmos w=1u l=1u
M6895 n3607 N528 VDD VDD pmos w=2u l=1u
M6896 n3607 N1 VDD VDD pmos w=2u l=1u
M6897 n3608 n3605 net2080 VSS nmos w=1u l=1u
M6898 net2080 n3609 VSS VSS nmos w=1u l=1u
M6899 n3608 n3605 VDD VDD pmos w=2u l=1u
M6900 n3608 n3609 VDD VDD pmos w=2u l=1u
M6901 n3605 n3611 net2081 VSS nmos w=1u l=1u
M6902 net2081 n3610 VSS VSS nmos w=1u l=1u
M6903 n3605 n3611 VDD VDD pmos w=2u l=1u
M6904 n3605 n3610 VDD VDD pmos w=2u l=1u
M6905 n3611 n3613 net2082 VSS nmos w=1u l=1u
M6906 net2082 n3612 VSS VSS nmos w=1u l=1u
M6907 n3611 n3613 VDD VDD pmos w=2u l=1u
M6908 n3611 n3612 VDD VDD pmos w=2u l=1u
M6909 net2083 n3451 VSS VSS nmos w=1u l=1u
M6910 net2084 n3452 VSS VSS nmos w=1u l=1u
M6911 n3610 net2085 VSS VSS nmos w=1u l=1u
M6912 net2085 n3451 net2086 VSS nmos w=1u l=1u
M6913 net2085 net2083 net2084 VSS nmos w=1u l=1u
M6914 net2086 net2084 VSS VSS nmos w=1u l=1u
M6915 net2085 net2083 net2087 VDD pmos w=2u l=1u
M6916 net2083 n3451 VDD VDD pmos w=2u l=1u
M6917 net2084 n3451 net2085 VDD pmos w=2u l=1u
M6918 net2084 n3452 VDD VDD pmos w=2u l=1u
M6919 n3610 net2085 VDD VDD pmos w=2u l=1u
M6920 net2087 net2084 VDD VDD pmos w=2u l=1u
M6921 n3609 n3615 net2088 VSS nmos w=1u l=1u
M6922 net2088 n3614 VSS VSS nmos w=1u l=1u
M6923 n3609 n3615 VDD VDD pmos w=2u l=1u
M6924 n3609 n3614 VDD VDD pmos w=2u l=1u
M6925 net2089 n3452 VSS VSS nmos w=1u l=1u
M6926 net2090 n3616 VSS VSS nmos w=1u l=1u
M6927 n3615 net2091 VSS VSS nmos w=1u l=1u
M6928 net2091 n3452 net2092 VSS nmos w=1u l=1u
M6929 net2091 net2089 net2090 VSS nmos w=1u l=1u
M6930 net2092 net2090 VSS VSS nmos w=1u l=1u
M6931 net2091 net2089 net2093 VDD pmos w=2u l=1u
M6932 net2089 n3452 VDD VDD pmos w=2u l=1u
M6933 net2090 n3452 net2091 VDD pmos w=2u l=1u
M6934 net2090 n3616 VDD VDD pmos w=2u l=1u
M6935 n3615 net2091 VDD VDD pmos w=2u l=1u
M6936 net2093 net2090 VDD VDD pmos w=2u l=1u
M6937 n3452 n2232 VSS VSS nmos w=1u l=1u
M6938 n3452 n3603 VSS VSS nmos w=1u l=1u
M6939 n3452 n2232 net2094 VDD pmos w=2u l=1u
M6940 net2094 n3603 VDD VDD pmos w=2u l=1u
M6941 n3616 n3451 VDD VDD pmos w=2u l=1u
M6942 n3616 n3451 VSS VSS nmos w=1u l=1u
M6943 n3451 n3450 net2095 VSS nmos w=1u l=1u
M6944 net2095 n3617 VSS VSS nmos w=1u l=1u
M6945 n3451 n3450 VDD VDD pmos w=2u l=1u
M6946 n3451 n3617 VDD VDD pmos w=2u l=1u
M6947 n3450 n3619 net2096 VSS nmos w=1u l=1u
M6948 net2096 n3618 VSS VSS nmos w=1u l=1u
M6949 n3450 n3619 VDD VDD pmos w=2u l=1u
M6950 n3450 n3618 VDD VDD pmos w=2u l=1u
M6951 n3619 n3621 net2097 VSS nmos w=1u l=1u
M6952 net2097 n3620 VSS VSS nmos w=1u l=1u
M6953 n3619 n3621 VDD VDD pmos w=2u l=1u
M6954 n3619 n3620 VDD VDD pmos w=2u l=1u
M6955 n3620 net2098 VSS VSS nmos w=1u l=1u
M6956 net2098 n3622 VSS VSS nmos w=1u l=1u
M6957 net2098 n3623 VSS VSS nmos w=1u l=1u
M6958 net2098 n3623 net2099 VDD pmos w=2u l=1u
M6959 n3620 net2098 VDD VDD pmos w=2u l=1u
M6960 net2099 n3622 VDD VDD pmos w=2u l=1u
M6961 net2100 n3462 VSS VSS nmos w=1u l=1u
M6962 net2101 n3463 VSS VSS nmos w=1u l=1u
M6963 n3618 net2102 VSS VSS nmos w=1u l=1u
M6964 net2102 n3462 net2103 VSS nmos w=1u l=1u
M6965 net2102 net2100 net2101 VSS nmos w=1u l=1u
M6966 net2103 net2101 VSS VSS nmos w=1u l=1u
M6967 net2102 net2100 net2104 VDD pmos w=2u l=1u
M6968 net2100 n3462 VDD VDD pmos w=2u l=1u
M6969 net2101 n3462 net2102 VDD pmos w=2u l=1u
M6970 net2101 n3463 VDD VDD pmos w=2u l=1u
M6971 n3618 net2102 VDD VDD pmos w=2u l=1u
M6972 net2104 net2101 VDD VDD pmos w=2u l=1u
M6973 n3617 n3625 net2105 VSS nmos w=1u l=1u
M6974 net2105 n3624 VSS VSS nmos w=1u l=1u
M6975 n3617 n3625 VDD VDD pmos w=2u l=1u
M6976 n3617 n3624 VDD VDD pmos w=2u l=1u
M6977 net2106 n3463 VSS VSS nmos w=1u l=1u
M6978 net2107 n3626 VSS VSS nmos w=1u l=1u
M6979 n3625 net2108 VSS VSS nmos w=1u l=1u
M6980 net2108 n3463 net2109 VSS nmos w=1u l=1u
M6981 net2108 net2106 net2107 VSS nmos w=1u l=1u
M6982 net2109 net2107 VSS VSS nmos w=1u l=1u
M6983 net2108 net2106 net2110 VDD pmos w=2u l=1u
M6984 net2106 n3463 VDD VDD pmos w=2u l=1u
M6985 net2107 n3463 net2108 VDD pmos w=2u l=1u
M6986 net2107 n3626 VDD VDD pmos w=2u l=1u
M6987 n3625 net2108 VDD VDD pmos w=2u l=1u
M6988 net2110 net2107 VDD VDD pmos w=2u l=1u
M6989 n3463 n2271 VSS VSS nmos w=1u l=1u
M6990 n3463 n3456 VSS VSS nmos w=1u l=1u
M6991 n3463 n2271 net2111 VDD pmos w=2u l=1u
M6992 net2111 n3456 VDD VDD pmos w=2u l=1u
M6993 n3626 n3462 VDD VDD pmos w=2u l=1u
M6994 n3626 n3462 VSS VSS nmos w=1u l=1u
M6995 n3462 n3461 net2112 VSS nmos w=1u l=1u
M6996 net2112 n3627 VSS VSS nmos w=1u l=1u
M6997 n3462 n3461 VDD VDD pmos w=2u l=1u
M6998 n3462 n3627 VDD VDD pmos w=2u l=1u
M6999 n3461 n3629 net2113 VSS nmos w=1u l=1u
M7000 net2113 n3628 VSS VSS nmos w=1u l=1u
M7001 n3461 n3629 VDD VDD pmos w=2u l=1u
M7002 n3461 n3628 VDD VDD pmos w=2u l=1u
M7003 n3629 n3631 net2114 VSS nmos w=1u l=1u
M7004 net2114 n3630 VSS VSS nmos w=1u l=1u
M7005 n3629 n3631 VDD VDD pmos w=2u l=1u
M7006 n3629 n3630 VDD VDD pmos w=2u l=1u
M7007 n3630 net2115 VSS VSS nmos w=1u l=1u
M7008 net2115 n3632 VSS VSS nmos w=1u l=1u
M7009 net2115 n3633 VSS VSS nmos w=1u l=1u
M7010 net2115 n3633 net2116 VDD pmos w=2u l=1u
M7011 n3630 net2115 VDD VDD pmos w=2u l=1u
M7012 net2116 n3632 VDD VDD pmos w=2u l=1u
M7013 net2117 n3472 VSS VSS nmos w=1u l=1u
M7014 net2118 n3473 VSS VSS nmos w=1u l=1u
M7015 n3628 net2119 VSS VSS nmos w=1u l=1u
M7016 net2119 n3472 net2120 VSS nmos w=1u l=1u
M7017 net2119 net2117 net2118 VSS nmos w=1u l=1u
M7018 net2120 net2118 VSS VSS nmos w=1u l=1u
M7019 net2119 net2117 net2121 VDD pmos w=2u l=1u
M7020 net2117 n3472 VDD VDD pmos w=2u l=1u
M7021 net2118 n3472 net2119 VDD pmos w=2u l=1u
M7022 net2118 n3473 VDD VDD pmos w=2u l=1u
M7023 n3628 net2119 VDD VDD pmos w=2u l=1u
M7024 net2121 net2118 VDD VDD pmos w=2u l=1u
M7025 n3473 n3634 VDD VDD pmos w=2u l=1u
M7026 n3473 n3634 VSS VSS nmos w=1u l=1u
M7027 n3627 n3636 net2122 VSS nmos w=1u l=1u
M7028 net2122 n3635 VSS VSS nmos w=1u l=1u
M7029 n3627 n3636 VDD VDD pmos w=2u l=1u
M7030 n3627 n3635 VDD VDD pmos w=2u l=1u
M7031 net2123 n3634 VSS VSS nmos w=1u l=1u
M7032 net2124 n3472 VSS VSS nmos w=1u l=1u
M7033 n3636 net2125 VSS VSS nmos w=1u l=1u
M7034 net2125 n3634 net2126 VSS nmos w=1u l=1u
M7035 net2125 net2123 net2124 VSS nmos w=1u l=1u
M7036 net2126 net2124 VSS VSS nmos w=1u l=1u
M7037 net2125 net2123 net2127 VDD pmos w=2u l=1u
M7038 net2123 n3634 VDD VDD pmos w=2u l=1u
M7039 net2124 n3634 net2125 VDD pmos w=2u l=1u
M7040 net2124 n3472 VDD VDD pmos w=2u l=1u
M7041 n3636 net2125 VDD VDD pmos w=2u l=1u
M7042 net2127 net2124 VDD VDD pmos w=2u l=1u
M7043 n3634 N477 net2128 VSS nmos w=1u l=1u
M7044 net2128 N52 VSS VSS nmos w=1u l=1u
M7045 n3634 N477 VDD VDD pmos w=2u l=1u
M7046 n3634 N52 VDD VDD pmos w=2u l=1u
M7047 n3472 n3471 net2129 VSS nmos w=1u l=1u
M7048 net2129 n3637 VSS VSS nmos w=1u l=1u
M7049 n3472 n3471 VDD VDD pmos w=2u l=1u
M7050 n3472 n3637 VDD VDD pmos w=2u l=1u
M7051 n3471 n3639 net2130 VSS nmos w=1u l=1u
M7052 net2130 n3638 VSS VSS nmos w=1u l=1u
M7053 n3471 n3639 VDD VDD pmos w=2u l=1u
M7054 n3471 n3638 VDD VDD pmos w=2u l=1u
M7055 n3639 n3641 net2131 VSS nmos w=1u l=1u
M7056 net2131 n3640 VSS VSS nmos w=1u l=1u
M7057 n3639 n3641 VDD VDD pmos w=2u l=1u
M7058 n3639 n3640 VDD VDD pmos w=2u l=1u
M7059 n3640 net2132 VSS VSS nmos w=1u l=1u
M7060 net2132 n3642 VSS VSS nmos w=1u l=1u
M7061 net2132 n3643 VSS VSS nmos w=1u l=1u
M7062 net2132 n3643 net2133 VDD pmos w=2u l=1u
M7063 n3640 net2132 VDD VDD pmos w=2u l=1u
M7064 net2133 n3642 VDD VDD pmos w=2u l=1u
M7065 net2134 n3482 VSS VSS nmos w=1u l=1u
M7066 net2135 n3483 VSS VSS nmos w=1u l=1u
M7067 n3638 net2136 VSS VSS nmos w=1u l=1u
M7068 net2136 n3482 net2137 VSS nmos w=1u l=1u
M7069 net2136 net2134 net2135 VSS nmos w=1u l=1u
M7070 net2137 net2135 VSS VSS nmos w=1u l=1u
M7071 net2136 net2134 net2138 VDD pmos w=2u l=1u
M7072 net2134 n3482 VDD VDD pmos w=2u l=1u
M7073 net2135 n3482 net2136 VDD pmos w=2u l=1u
M7074 net2135 n3483 VDD VDD pmos w=2u l=1u
M7075 n3638 net2136 VDD VDD pmos w=2u l=1u
M7076 net2138 net2135 VDD VDD pmos w=2u l=1u
M7077 n3483 n3644 VDD VDD pmos w=2u l=1u
M7078 n3483 n3644 VSS VSS nmos w=1u l=1u
M7079 n3637 n3646 net2139 VSS nmos w=1u l=1u
M7080 net2139 n3645 VSS VSS nmos w=1u l=1u
M7081 n3637 n3646 VDD VDD pmos w=2u l=1u
M7082 n3637 n3645 VDD VDD pmos w=2u l=1u
M7083 net2140 n3644 VSS VSS nmos w=1u l=1u
M7084 net2141 n3482 VSS VSS nmos w=1u l=1u
M7085 n3646 net2142 VSS VSS nmos w=1u l=1u
M7086 net2142 n3644 net2143 VSS nmos w=1u l=1u
M7087 net2142 net2140 net2141 VSS nmos w=1u l=1u
M7088 net2143 net2141 VSS VSS nmos w=1u l=1u
M7089 net2142 net2140 net2144 VDD pmos w=2u l=1u
M7090 net2140 n3644 VDD VDD pmos w=2u l=1u
M7091 net2141 n3644 net2142 VDD pmos w=2u l=1u
M7092 net2141 n3482 VDD VDD pmos w=2u l=1u
M7093 n3646 net2142 VDD VDD pmos w=2u l=1u
M7094 net2144 net2141 VDD VDD pmos w=2u l=1u
M7095 n3644 N460 net2145 VSS nmos w=1u l=1u
M7096 net2145 N69 VSS VSS nmos w=1u l=1u
M7097 n3644 N460 VDD VDD pmos w=2u l=1u
M7098 n3644 N69 VDD VDD pmos w=2u l=1u
M7099 n3482 n3481 net2146 VSS nmos w=1u l=1u
M7100 net2146 n3647 VSS VSS nmos w=1u l=1u
M7101 n3482 n3481 VDD VDD pmos w=2u l=1u
M7102 n3482 n3647 VDD VDD pmos w=2u l=1u
M7103 n3481 n3649 net2147 VSS nmos w=1u l=1u
M7104 net2147 n3648 VSS VSS nmos w=1u l=1u
M7105 n3481 n3649 VDD VDD pmos w=2u l=1u
M7106 n3481 n3648 VDD VDD pmos w=2u l=1u
M7107 n3649 n3651 net2148 VSS nmos w=1u l=1u
M7108 net2148 n3650 VSS VSS nmos w=1u l=1u
M7109 n3649 n3651 VDD VDD pmos w=2u l=1u
M7110 n3649 n3650 VDD VDD pmos w=2u l=1u
M7111 n3650 net2149 VSS VSS nmos w=1u l=1u
M7112 net2149 n3652 VSS VSS nmos w=1u l=1u
M7113 net2149 n3653 VSS VSS nmos w=1u l=1u
M7114 net2149 n3653 net2150 VDD pmos w=2u l=1u
M7115 n3650 net2149 VDD VDD pmos w=2u l=1u
M7116 net2150 n3652 VDD VDD pmos w=2u l=1u
M7117 net2151 n3492 VSS VSS nmos w=1u l=1u
M7118 net2152 n3493 VSS VSS nmos w=1u l=1u
M7119 n3648 net2153 VSS VSS nmos w=1u l=1u
M7120 net2153 n3492 net2154 VSS nmos w=1u l=1u
M7121 net2153 net2151 net2152 VSS nmos w=1u l=1u
M7122 net2154 net2152 VSS VSS nmos w=1u l=1u
M7123 net2153 net2151 net2155 VDD pmos w=2u l=1u
M7124 net2151 n3492 VDD VDD pmos w=2u l=1u
M7125 net2152 n3492 net2153 VDD pmos w=2u l=1u
M7126 net2152 n3493 VDD VDD pmos w=2u l=1u
M7127 n3648 net2153 VDD VDD pmos w=2u l=1u
M7128 net2155 net2152 VDD VDD pmos w=2u l=1u
M7129 n3493 n3654 VDD VDD pmos w=2u l=1u
M7130 n3493 n3654 VSS VSS nmos w=1u l=1u
M7131 n3647 n3656 net2156 VSS nmos w=1u l=1u
M7132 net2156 n3655 VSS VSS nmos w=1u l=1u
M7133 n3647 n3656 VDD VDD pmos w=2u l=1u
M7134 n3647 n3655 VDD VDD pmos w=2u l=1u
M7135 net2157 n3654 VSS VSS nmos w=1u l=1u
M7136 net2158 n3492 VSS VSS nmos w=1u l=1u
M7137 n3656 net2159 VSS VSS nmos w=1u l=1u
M7138 net2159 n3654 net2160 VSS nmos w=1u l=1u
M7139 net2159 net2157 net2158 VSS nmos w=1u l=1u
M7140 net2160 net2158 VSS VSS nmos w=1u l=1u
M7141 net2159 net2157 net2161 VDD pmos w=2u l=1u
M7142 net2157 n3654 VDD VDD pmos w=2u l=1u
M7143 net2158 n3654 net2159 VDD pmos w=2u l=1u
M7144 net2158 n3492 VDD VDD pmos w=2u l=1u
M7145 n3656 net2159 VDD VDD pmos w=2u l=1u
M7146 net2161 net2158 VDD VDD pmos w=2u l=1u
M7147 n3654 N443 net2162 VSS nmos w=1u l=1u
M7148 net2162 N86 VSS VSS nmos w=1u l=1u
M7149 n3654 N443 VDD VDD pmos w=2u l=1u
M7150 n3654 N86 VDD VDD pmos w=2u l=1u
M7151 n3492 n3491 net2163 VSS nmos w=1u l=1u
M7152 net2163 n3657 VSS VSS nmos w=1u l=1u
M7153 n3492 n3491 VDD VDD pmos w=2u l=1u
M7154 n3492 n3657 VDD VDD pmos w=2u l=1u
M7155 n3491 n3659 net2164 VSS nmos w=1u l=1u
M7156 net2164 n3658 VSS VSS nmos w=1u l=1u
M7157 n3491 n3659 VDD VDD pmos w=2u l=1u
M7158 n3491 n3658 VDD VDD pmos w=2u l=1u
M7159 n3659 n3661 net2165 VSS nmos w=1u l=1u
M7160 net2165 n3660 VSS VSS nmos w=1u l=1u
M7161 n3659 n3661 VDD VDD pmos w=2u l=1u
M7162 n3659 n3660 VDD VDD pmos w=2u l=1u
M7163 n3660 net2166 VSS VSS nmos w=1u l=1u
M7164 net2166 n3662 VSS VSS nmos w=1u l=1u
M7165 net2166 n3663 VSS VSS nmos w=1u l=1u
M7166 net2166 n3663 net2167 VDD pmos w=2u l=1u
M7167 n3660 net2166 VDD VDD pmos w=2u l=1u
M7168 net2167 n3662 VDD VDD pmos w=2u l=1u
M7169 net2168 n3502 VSS VSS nmos w=1u l=1u
M7170 net2169 n3503 VSS VSS nmos w=1u l=1u
M7171 n3658 net2170 VSS VSS nmos w=1u l=1u
M7172 net2170 n3502 net2171 VSS nmos w=1u l=1u
M7173 net2170 net2168 net2169 VSS nmos w=1u l=1u
M7174 net2171 net2169 VSS VSS nmos w=1u l=1u
M7175 net2170 net2168 net2172 VDD pmos w=2u l=1u
M7176 net2168 n3502 VDD VDD pmos w=2u l=1u
M7177 net2169 n3502 net2170 VDD pmos w=2u l=1u
M7178 net2169 n3503 VDD VDD pmos w=2u l=1u
M7179 n3658 net2170 VDD VDD pmos w=2u l=1u
M7180 net2172 net2169 VDD VDD pmos w=2u l=1u
M7181 n3503 n3664 VDD VDD pmos w=2u l=1u
M7182 n3503 n3664 VSS VSS nmos w=1u l=1u
M7183 n3657 n3666 net2173 VSS nmos w=1u l=1u
M7184 net2173 n3665 VSS VSS nmos w=1u l=1u
M7185 n3657 n3666 VDD VDD pmos w=2u l=1u
M7186 n3657 n3665 VDD VDD pmos w=2u l=1u
M7187 net2174 n3664 VSS VSS nmos w=1u l=1u
M7188 net2175 n3502 VSS VSS nmos w=1u l=1u
M7189 n3666 net2176 VSS VSS nmos w=1u l=1u
M7190 net2176 n3664 net2177 VSS nmos w=1u l=1u
M7191 net2176 net2174 net2175 VSS nmos w=1u l=1u
M7192 net2177 net2175 VSS VSS nmos w=1u l=1u
M7193 net2176 net2174 net2178 VDD pmos w=2u l=1u
M7194 net2174 n3664 VDD VDD pmos w=2u l=1u
M7195 net2175 n3664 net2176 VDD pmos w=2u l=1u
M7196 net2175 n3502 VDD VDD pmos w=2u l=1u
M7197 n3666 net2176 VDD VDD pmos w=2u l=1u
M7198 net2178 net2175 VDD VDD pmos w=2u l=1u
M7199 n3664 N426 net2179 VSS nmos w=1u l=1u
M7200 net2179 N103 VSS VSS nmos w=1u l=1u
M7201 n3664 N426 VDD VDD pmos w=2u l=1u
M7202 n3664 N103 VDD VDD pmos w=2u l=1u
M7203 n3502 n3501 net2180 VSS nmos w=1u l=1u
M7204 net2180 n3667 VSS VSS nmos w=1u l=1u
M7205 n3502 n3501 VDD VDD pmos w=2u l=1u
M7206 n3502 n3667 VDD VDD pmos w=2u l=1u
M7207 n3501 n3669 net2181 VSS nmos w=1u l=1u
M7208 net2181 n3668 VSS VSS nmos w=1u l=1u
M7209 n3501 n3669 VDD VDD pmos w=2u l=1u
M7210 n3501 n3668 VDD VDD pmos w=2u l=1u
M7211 n3669 n3671 net2182 VSS nmos w=1u l=1u
M7212 net2182 n3670 VSS VSS nmos w=1u l=1u
M7213 n3669 n3671 VDD VDD pmos w=2u l=1u
M7214 n3669 n3670 VDD VDD pmos w=2u l=1u
M7215 n3670 net2183 VSS VSS nmos w=1u l=1u
M7216 net2183 n3672 VSS VSS nmos w=1u l=1u
M7217 net2183 n3673 VSS VSS nmos w=1u l=1u
M7218 net2183 n3673 net2184 VDD pmos w=2u l=1u
M7219 n3670 net2183 VDD VDD pmos w=2u l=1u
M7220 net2184 n3672 VDD VDD pmos w=2u l=1u
M7221 net2185 n3512 VSS VSS nmos w=1u l=1u
M7222 net2186 n3513 VSS VSS nmos w=1u l=1u
M7223 n3668 net2187 VSS VSS nmos w=1u l=1u
M7224 net2187 n3512 net2188 VSS nmos w=1u l=1u
M7225 net2187 net2185 net2186 VSS nmos w=1u l=1u
M7226 net2188 net2186 VSS VSS nmos w=1u l=1u
M7227 net2187 net2185 net2189 VDD pmos w=2u l=1u
M7228 net2185 n3512 VDD VDD pmos w=2u l=1u
M7229 net2186 n3512 net2187 VDD pmos w=2u l=1u
M7230 net2186 n3513 VDD VDD pmos w=2u l=1u
M7231 n3668 net2187 VDD VDD pmos w=2u l=1u
M7232 net2189 net2186 VDD VDD pmos w=2u l=1u
M7233 n3513 n3674 VDD VDD pmos w=2u l=1u
M7234 n3513 n3674 VSS VSS nmos w=1u l=1u
M7235 n3667 n3676 net2190 VSS nmos w=1u l=1u
M7236 net2190 n3675 VSS VSS nmos w=1u l=1u
M7237 n3667 n3676 VDD VDD pmos w=2u l=1u
M7238 n3667 n3675 VDD VDD pmos w=2u l=1u
M7239 net2191 n3674 VSS VSS nmos w=1u l=1u
M7240 net2192 n3512 VSS VSS nmos w=1u l=1u
M7241 n3676 net2193 VSS VSS nmos w=1u l=1u
M7242 net2193 n3674 net2194 VSS nmos w=1u l=1u
M7243 net2193 net2191 net2192 VSS nmos w=1u l=1u
M7244 net2194 net2192 VSS VSS nmos w=1u l=1u
M7245 net2193 net2191 net2195 VDD pmos w=2u l=1u
M7246 net2191 n3674 VDD VDD pmos w=2u l=1u
M7247 net2192 n3674 net2193 VDD pmos w=2u l=1u
M7248 net2192 n3512 VDD VDD pmos w=2u l=1u
M7249 n3676 net2193 VDD VDD pmos w=2u l=1u
M7250 net2195 net2192 VDD VDD pmos w=2u l=1u
M7251 n3674 N409 net2196 VSS nmos w=1u l=1u
M7252 net2196 N120 VSS VSS nmos w=1u l=1u
M7253 n3674 N409 VDD VDD pmos w=2u l=1u
M7254 n3674 N120 VDD VDD pmos w=2u l=1u
M7255 n3512 n3511 net2197 VSS nmos w=1u l=1u
M7256 net2197 n3677 VSS VSS nmos w=1u l=1u
M7257 n3512 n3511 VDD VDD pmos w=2u l=1u
M7258 n3512 n3677 VDD VDD pmos w=2u l=1u
M7259 n3511 n3679 net2198 VSS nmos w=1u l=1u
M7260 net2198 n3678 VSS VSS nmos w=1u l=1u
M7261 n3511 n3679 VDD VDD pmos w=2u l=1u
M7262 n3511 n3678 VDD VDD pmos w=2u l=1u
M7263 n3679 n3681 net2199 VSS nmos w=1u l=1u
M7264 net2199 n3680 VSS VSS nmos w=1u l=1u
M7265 n3679 n3681 VDD VDD pmos w=2u l=1u
M7266 n3679 n3680 VDD VDD pmos w=2u l=1u
M7267 n3680 net2200 VSS VSS nmos w=1u l=1u
M7268 net2200 n3682 VSS VSS nmos w=1u l=1u
M7269 net2200 n3683 VSS VSS nmos w=1u l=1u
M7270 net2200 n3683 net2201 VDD pmos w=2u l=1u
M7271 n3680 net2200 VDD VDD pmos w=2u l=1u
M7272 net2201 n3682 VDD VDD pmos w=2u l=1u
M7273 net2202 n3522 VSS VSS nmos w=1u l=1u
M7274 net2203 n3523 VSS VSS nmos w=1u l=1u
M7275 n3678 net2204 VSS VSS nmos w=1u l=1u
M7276 net2204 n3522 net2205 VSS nmos w=1u l=1u
M7277 net2204 net2202 net2203 VSS nmos w=1u l=1u
M7278 net2205 net2203 VSS VSS nmos w=1u l=1u
M7279 net2204 net2202 net2206 VDD pmos w=2u l=1u
M7280 net2202 n3522 VDD VDD pmos w=2u l=1u
M7281 net2203 n3522 net2204 VDD pmos w=2u l=1u
M7282 net2203 n3523 VDD VDD pmos w=2u l=1u
M7283 n3678 net2204 VDD VDD pmos w=2u l=1u
M7284 net2206 net2203 VDD VDD pmos w=2u l=1u
M7285 n3523 n3684 VDD VDD pmos w=2u l=1u
M7286 n3523 n3684 VSS VSS nmos w=1u l=1u
M7287 n3677 n3686 net2207 VSS nmos w=1u l=1u
M7288 net2207 n3685 VSS VSS nmos w=1u l=1u
M7289 n3677 n3686 VDD VDD pmos w=2u l=1u
M7290 n3677 n3685 VDD VDD pmos w=2u l=1u
M7291 net2208 n3684 VSS VSS nmos w=1u l=1u
M7292 net2209 n3522 VSS VSS nmos w=1u l=1u
M7293 n3686 net2210 VSS VSS nmos w=1u l=1u
M7294 net2210 n3684 net2211 VSS nmos w=1u l=1u
M7295 net2210 net2208 net2209 VSS nmos w=1u l=1u
M7296 net2211 net2209 VSS VSS nmos w=1u l=1u
M7297 net2210 net2208 net2212 VDD pmos w=2u l=1u
M7298 net2208 n3684 VDD VDD pmos w=2u l=1u
M7299 net2209 n3684 net2210 VDD pmos w=2u l=1u
M7300 net2209 n3522 VDD VDD pmos w=2u l=1u
M7301 n3686 net2210 VDD VDD pmos w=2u l=1u
M7302 net2212 net2209 VDD VDD pmos w=2u l=1u
M7303 n3684 N392 net2213 VSS nmos w=1u l=1u
M7304 net2213 N137 VSS VSS nmos w=1u l=1u
M7305 n3684 N392 VDD VDD pmos w=2u l=1u
M7306 n3684 N137 VDD VDD pmos w=2u l=1u
M7307 n3522 n3521 net2214 VSS nmos w=1u l=1u
M7308 net2214 n3687 VSS VSS nmos w=1u l=1u
M7309 n3522 n3521 VDD VDD pmos w=2u l=1u
M7310 n3522 n3687 VDD VDD pmos w=2u l=1u
M7311 n3521 n3689 net2215 VSS nmos w=1u l=1u
M7312 net2215 n3688 VSS VSS nmos w=1u l=1u
M7313 n3521 n3689 VDD VDD pmos w=2u l=1u
M7314 n3521 n3688 VDD VDD pmos w=2u l=1u
M7315 n3689 n3691 net2216 VSS nmos w=1u l=1u
M7316 net2216 n3690 VSS VSS nmos w=1u l=1u
M7317 n3689 n3691 VDD VDD pmos w=2u l=1u
M7318 n3689 n3690 VDD VDD pmos w=2u l=1u
M7319 n3690 net2217 VSS VSS nmos w=1u l=1u
M7320 net2217 n3692 VSS VSS nmos w=1u l=1u
M7321 net2217 n3693 VSS VSS nmos w=1u l=1u
M7322 net2217 n3693 net2218 VDD pmos w=2u l=1u
M7323 n3690 net2217 VDD VDD pmos w=2u l=1u
M7324 net2218 n3692 VDD VDD pmos w=2u l=1u
M7325 net2219 n3532 VSS VSS nmos w=1u l=1u
M7326 net2220 n3533 VSS VSS nmos w=1u l=1u
M7327 n3688 net2221 VSS VSS nmos w=1u l=1u
M7328 net2221 n3532 net2222 VSS nmos w=1u l=1u
M7329 net2221 net2219 net2220 VSS nmos w=1u l=1u
M7330 net2222 net2220 VSS VSS nmos w=1u l=1u
M7331 net2221 net2219 net2223 VDD pmos w=2u l=1u
M7332 net2219 n3532 VDD VDD pmos w=2u l=1u
M7333 net2220 n3532 net2221 VDD pmos w=2u l=1u
M7334 net2220 n3533 VDD VDD pmos w=2u l=1u
M7335 n3688 net2221 VDD VDD pmos w=2u l=1u
M7336 net2223 net2220 VDD VDD pmos w=2u l=1u
M7337 n3532 n3694 VDD VDD pmos w=2u l=1u
M7338 n3532 n3694 VSS VSS nmos w=1u l=1u
M7339 n3687 n3696 net2224 VSS nmos w=1u l=1u
M7340 net2224 n3695 VSS VSS nmos w=1u l=1u
M7341 n3687 n3696 VDD VDD pmos w=2u l=1u
M7342 n3687 n3695 VDD VDD pmos w=2u l=1u
M7343 net2225 n3533 VSS VSS nmos w=1u l=1u
M7344 net2226 n3694 VSS VSS nmos w=1u l=1u
M7345 n3696 net2227 VSS VSS nmos w=1u l=1u
M7346 net2227 n3533 net2228 VSS nmos w=1u l=1u
M7347 net2227 net2225 net2226 VSS nmos w=1u l=1u
M7348 net2228 net2226 VSS VSS nmos w=1u l=1u
M7349 net2227 net2225 net2229 VDD pmos w=2u l=1u
M7350 net2225 n3533 VDD VDD pmos w=2u l=1u
M7351 net2226 n3533 net2227 VDD pmos w=2u l=1u
M7352 net2226 n3694 VDD VDD pmos w=2u l=1u
M7353 n3696 net2227 VDD VDD pmos w=2u l=1u
M7354 net2229 net2226 VDD VDD pmos w=2u l=1u
M7355 n3533 N375 net2230 VSS nmos w=1u l=1u
M7356 net2230 N154 VSS VSS nmos w=1u l=1u
M7357 n3533 N375 VDD VDD pmos w=2u l=1u
M7358 n3533 N154 VDD VDD pmos w=2u l=1u
M7359 n3694 n3531 net2231 VSS nmos w=1u l=1u
M7360 net2231 n3697 VSS VSS nmos w=1u l=1u
M7361 n3694 n3531 VDD VDD pmos w=2u l=1u
M7362 n3694 n3697 VDD VDD pmos w=2u l=1u
M7363 n3531 n3699 net2232 VSS nmos w=1u l=1u
M7364 net2232 n3698 VSS VSS nmos w=1u l=1u
M7365 n3531 n3699 VDD VDD pmos w=2u l=1u
M7366 n3531 n3698 VDD VDD pmos w=2u l=1u
M7367 n3699 n3701 net2233 VSS nmos w=1u l=1u
M7368 net2233 n3700 VSS VSS nmos w=1u l=1u
M7369 n3699 n3701 VDD VDD pmos w=2u l=1u
M7370 n3699 n3700 VDD VDD pmos w=2u l=1u
M7371 n3700 net2234 VSS VSS nmos w=1u l=1u
M7372 net2234 n3702 VSS VSS nmos w=1u l=1u
M7373 net2234 n3703 VSS VSS nmos w=1u l=1u
M7374 net2234 n3703 net2235 VDD pmos w=2u l=1u
M7375 n3700 net2234 VDD VDD pmos w=2u l=1u
M7376 net2235 n3702 VDD VDD pmos w=2u l=1u
M7377 net2236 n3542 VSS VSS nmos w=1u l=1u
M7378 net2237 n3543 VSS VSS nmos w=1u l=1u
M7379 n3698 net2238 VSS VSS nmos w=1u l=1u
M7380 net2238 n3542 net2239 VSS nmos w=1u l=1u
M7381 net2238 net2236 net2237 VSS nmos w=1u l=1u
M7382 net2239 net2237 VSS VSS nmos w=1u l=1u
M7383 net2238 net2236 net2240 VDD pmos w=2u l=1u
M7384 net2236 n3542 VDD VDD pmos w=2u l=1u
M7385 net2237 n3542 net2238 VDD pmos w=2u l=1u
M7386 net2237 n3543 VDD VDD pmos w=2u l=1u
M7387 n3698 net2238 VDD VDD pmos w=2u l=1u
M7388 net2240 net2237 VDD VDD pmos w=2u l=1u
M7389 n3543 n3704 VDD VDD pmos w=2u l=1u
M7390 n3543 n3704 VSS VSS nmos w=1u l=1u
M7391 n3697 n3706 net2241 VSS nmos w=1u l=1u
M7392 net2241 n3705 VSS VSS nmos w=1u l=1u
M7393 n3697 n3706 VDD VDD pmos w=2u l=1u
M7394 n3697 n3705 VDD VDD pmos w=2u l=1u
M7395 net2242 n3704 VSS VSS nmos w=1u l=1u
M7396 net2243 n3542 VSS VSS nmos w=1u l=1u
M7397 n3706 net2244 VSS VSS nmos w=1u l=1u
M7398 net2244 n3704 net2245 VSS nmos w=1u l=1u
M7399 net2244 net2242 net2243 VSS nmos w=1u l=1u
M7400 net2245 net2243 VSS VSS nmos w=1u l=1u
M7401 net2244 net2242 net2246 VDD pmos w=2u l=1u
M7402 net2242 n3704 VDD VDD pmos w=2u l=1u
M7403 net2243 n3704 net2244 VDD pmos w=2u l=1u
M7404 net2243 n3542 VDD VDD pmos w=2u l=1u
M7405 n3706 net2244 VDD VDD pmos w=2u l=1u
M7406 net2246 net2243 VDD VDD pmos w=2u l=1u
M7407 n3704 N358 net2247 VSS nmos w=1u l=1u
M7408 net2247 N171 VSS VSS nmos w=1u l=1u
M7409 n3704 N358 VDD VDD pmos w=2u l=1u
M7410 n3704 N171 VDD VDD pmos w=2u l=1u
M7411 n3542 n3541 net2248 VSS nmos w=1u l=1u
M7412 net2248 n3707 VSS VSS nmos w=1u l=1u
M7413 n3542 n3541 VDD VDD pmos w=2u l=1u
M7414 n3542 n3707 VDD VDD pmos w=2u l=1u
M7415 n3541 n3709 net2249 VSS nmos w=1u l=1u
M7416 net2249 n3708 VSS VSS nmos w=1u l=1u
M7417 n3541 n3709 VDD VDD pmos w=2u l=1u
M7418 n3541 n3708 VDD VDD pmos w=2u l=1u
M7419 n3709 n3711 net2250 VSS nmos w=1u l=1u
M7420 net2250 n3710 VSS VSS nmos w=1u l=1u
M7421 n3709 n3711 VDD VDD pmos w=2u l=1u
M7422 n3709 n3710 VDD VDD pmos w=2u l=1u
M7423 n3710 n3713 net2251 VSS nmos w=1u l=1u
M7424 net2251 n3712 VSS VSS nmos w=1u l=1u
M7425 n3710 n3713 VDD VDD pmos w=2u l=1u
M7426 n3710 n3712 VDD VDD pmos w=2u l=1u
M7427 net2252 n3552 VSS VSS nmos w=1u l=1u
M7428 net2253 n3553 VSS VSS nmos w=1u l=1u
M7429 n3708 net2254 VSS VSS nmos w=1u l=1u
M7430 net2254 n3552 net2255 VSS nmos w=1u l=1u
M7431 net2254 net2252 net2253 VSS nmos w=1u l=1u
M7432 net2255 net2253 VSS VSS nmos w=1u l=1u
M7433 net2254 net2252 net2256 VDD pmos w=2u l=1u
M7434 net2252 n3552 VDD VDD pmos w=2u l=1u
M7435 net2253 n3552 net2254 VDD pmos w=2u l=1u
M7436 net2253 n3553 VDD VDD pmos w=2u l=1u
M7437 n3708 net2254 VDD VDD pmos w=2u l=1u
M7438 net2256 net2253 VDD VDD pmos w=2u l=1u
M7439 n3553 n3714 VDD VDD pmos w=2u l=1u
M7440 n3553 n3714 VSS VSS nmos w=1u l=1u
M7441 n3707 n3716 net2257 VSS nmos w=1u l=1u
M7442 net2257 n3715 VSS VSS nmos w=1u l=1u
M7443 n3707 n3716 VDD VDD pmos w=2u l=1u
M7444 n3707 n3715 VDD VDD pmos w=2u l=1u
M7445 net2258 n3714 VSS VSS nmos w=1u l=1u
M7446 net2259 n3552 VSS VSS nmos w=1u l=1u
M7447 n3716 net2260 VSS VSS nmos w=1u l=1u
M7448 net2260 n3714 net2261 VSS nmos w=1u l=1u
M7449 net2260 net2258 net2259 VSS nmos w=1u l=1u
M7450 net2261 net2259 VSS VSS nmos w=1u l=1u
M7451 net2260 net2258 net2262 VDD pmos w=2u l=1u
M7452 net2258 n3714 VDD VDD pmos w=2u l=1u
M7453 net2259 n3714 net2260 VDD pmos w=2u l=1u
M7454 net2259 n3552 VDD VDD pmos w=2u l=1u
M7455 n3716 net2260 VDD VDD pmos w=2u l=1u
M7456 net2262 net2259 VDD VDD pmos w=2u l=1u
M7457 n3714 N341 net2263 VSS nmos w=1u l=1u
M7458 net2263 N188 VSS VSS nmos w=1u l=1u
M7459 n3714 N341 VDD VDD pmos w=2u l=1u
M7460 n3714 N188 VDD VDD pmos w=2u l=1u
M7461 n3552 n3551 net2264 VSS nmos w=1u l=1u
M7462 net2264 n3717 VSS VSS nmos w=1u l=1u
M7463 n3552 n3551 VDD VDD pmos w=2u l=1u
M7464 n3552 n3717 VDD VDD pmos w=2u l=1u
M7465 n3551 n3719 net2265 VSS nmos w=1u l=1u
M7466 net2265 n3718 VSS VSS nmos w=1u l=1u
M7467 n3551 n3719 VDD VDD pmos w=2u l=1u
M7468 n3551 n3718 VDD VDD pmos w=2u l=1u
M7469 n3719 net2266 VSS VSS nmos w=1u l=1u
M7470 net2266 n3720 VSS VSS nmos w=1u l=1u
M7471 net2266 n3721 VSS VSS nmos w=1u l=1u
M7472 net2266 n3721 net2267 VDD pmos w=2u l=1u
M7473 n3719 net2266 VDD VDD pmos w=2u l=1u
M7474 net2267 n3720 VDD VDD pmos w=2u l=1u
M7475 n3718 net2268 VSS VSS nmos w=1u l=1u
M7476 net2269 n3722 VSS VSS nmos w=1u l=1u
M7477 net2268 n3580 net2269 VSS nmos w=1u l=1u
M7478 net2268 n3722 VDD VDD pmos w=2u l=1u
M7479 net2268 n3580 VDD VDD pmos w=2u l=1u
M7480 n3718 net2268 VDD VDD pmos w=2u l=1u
M7481 n3717 n3724 net2270 VSS nmos w=1u l=1u
M7482 net2270 n3723 VSS VSS nmos w=1u l=1u
M7483 n3717 n3724 VDD VDD pmos w=2u l=1u
M7484 n3717 n3723 VDD VDD pmos w=2u l=1u
M7485 n3724 n3580 net2271 VSS nmos w=1u l=1u
M7486 net2271 n3722 VSS VSS nmos w=1u l=1u
M7487 n3724 n3580 VDD VDD pmos w=2u l=1u
M7488 n3724 n3722 VDD VDD pmos w=2u l=1u
M7489 n3580 n3726 net2272 VSS nmos w=1u l=1u
M7490 net2272 n3725 VSS VSS nmos w=1u l=1u
M7491 n3580 n3726 VDD VDD pmos w=2u l=1u
M7492 n3580 n3725 VDD VDD pmos w=2u l=1u
M7493 n3726 N324 net2273 VSS nmos w=1u l=1u
M7494 net2273 N205 VSS VSS nmos w=1u l=1u
M7495 n3726 N324 VDD VDD pmos w=2u l=1u
M7496 n3726 N205 VDD VDD pmos w=2u l=1u
M7497 n3722 N205 net2274 VSS nmos w=1u l=1u
M7498 net2274 n3727 VSS VSS nmos w=1u l=1u
M7499 n3722 N205 VDD VDD pmos w=2u l=1u
M7500 n3722 n3727 VDD VDD pmos w=2u l=1u
M7501 n3727 n3257 VSS VSS nmos w=1u l=1u
M7502 n3727 n3725 VSS VSS nmos w=1u l=1u
M7503 n3727 n3257 net2275 VDD pmos w=2u l=1u
M7504 net2275 n3725 VDD VDD pmos w=2u l=1u
M7505 n3725 n3561 VSS VSS nmos w=1u l=1u
M7506 n3725 n3728 VSS VSS nmos w=1u l=1u
M7507 n3725 n3561 net2276 VDD pmos w=2u l=1u
M7508 net2276 n3728 VDD VDD pmos w=2u l=1u
M7509 n3561 n3730 VSS VSS nmos w=1u l=1u
M7510 n3561 n3729 VSS VSS nmos w=1u l=1u
M7511 n3561 n3730 net2277 VDD pmos w=2u l=1u
M7512 net2277 n3729 VDD VDD pmos w=2u l=1u
M7513 n3728 net2278 VSS VSS nmos w=1u l=1u
M7514 net2279 n3729 VSS VSS nmos w=1u l=1u
M7515 net2278 n3730 net2279 VSS nmos w=1u l=1u
M7516 net2278 n3729 VDD VDD pmos w=2u l=1u
M7517 net2278 n3730 VDD VDD pmos w=2u l=1u
M7518 n3728 net2278 VDD VDD pmos w=2u l=1u
M7519 n3729 n3731 net2280 VSS nmos w=1u l=1u
M7520 net2280 n3578 VSS VSS nmos w=1u l=1u
M7521 n3729 n3731 VDD VDD pmos w=2u l=1u
M7522 n3729 n3578 VDD VDD pmos w=2u l=1u
M7523 n3731 N222 net2281 VSS nmos w=1u l=1u
M7524 net2281 n3732 VSS VSS nmos w=1u l=1u
M7525 n3731 N222 VDD VDD pmos w=2u l=1u
M7526 n3731 n3732 VDD VDD pmos w=2u l=1u
M7527 n3732 n3411 VSS VSS nmos w=1u l=1u
M7528 n3732 n3733 VSS VSS nmos w=1u l=1u
M7529 n3732 n3411 net2282 VDD pmos w=2u l=1u
M7530 net2282 n3733 VDD VDD pmos w=2u l=1u
M7531 n3578 n3734 net2283 VSS nmos w=1u l=1u
M7532 net2283 n3733 VSS VSS nmos w=1u l=1u
M7533 n3578 n3734 VDD VDD pmos w=2u l=1u
M7534 n3578 n3733 VDD VDD pmos w=2u l=1u
M7535 n3734 N307 net2284 VSS nmos w=1u l=1u
M7536 net2284 N222 VSS VSS nmos w=1u l=1u
M7537 n3734 N307 VDD VDD pmos w=2u l=1u
M7538 n3734 N222 VDD VDD pmos w=2u l=1u
M7539 n3733 net2285 VSS VSS nmos w=1u l=1u
M7540 net2286 n3735 VSS VSS nmos w=1u l=1u
M7541 net2285 n3579 net2286 VSS nmos w=1u l=1u
M7542 net2285 n3735 VDD VDD pmos w=2u l=1u
M7543 net2285 n3579 VDD VDD pmos w=2u l=1u
M7544 n3733 net2285 VDD VDD pmos w=2u l=1u
M7545 n3735 n3737 net2287 VSS nmos w=1u l=1u
M7546 net2287 n3736 VSS VSS nmos w=1u l=1u
M7547 n3735 n3737 VDD VDD pmos w=2u l=1u
M7548 n3735 n3736 VDD VDD pmos w=2u l=1u
M7549 n3579 n3739 net2288 VSS nmos w=1u l=1u
M7550 net2288 n3738 VSS VSS nmos w=1u l=1u
M7551 n3579 n3739 VDD VDD pmos w=2u l=1u
M7552 n3579 n3738 VDD VDD pmos w=2u l=1u
M7553 n3739 N239 net2289 VSS nmos w=1u l=1u
M7554 net2289 n3576 VSS VSS nmos w=1u l=1u
M7555 n3739 N239 VDD VDD pmos w=2u l=1u
M7556 n3739 n3576 VDD VDD pmos w=2u l=1u
M7557 n3576 n3574 VDD VDD pmos w=2u l=1u
M7558 n3576 n3574 VSS VSS nmos w=1u l=1u
M7559 n3574 n3737 net2290 VSS nmos w=1u l=1u
M7560 net2290 N290 VSS VSS nmos w=1u l=1u
M7561 n3574 n3737 VDD VDD pmos w=2u l=1u
M7562 n3574 N290 VDD VDD pmos w=2u l=1u
M7563 n3737 n3741 net2291 VSS nmos w=1u l=1u
M7564 net2291 n3740 VSS VSS nmos w=1u l=1u
M7565 n3737 n3741 VDD VDD pmos w=2u l=1u
M7566 n3737 n3740 VDD VDD pmos w=2u l=1u
M7567 n3740 n2275 VSS VSS nmos w=1u l=1u
M7568 n3740 n2228 VSS VSS nmos w=1u l=1u
M7569 n3740 n2275 net2292 VDD pmos w=2u l=1u
M7570 net2292 n2228 VDD VDD pmos w=2u l=1u
M7571 n3738 n3742 VSS VSS nmos w=1u l=1u
M7572 n3738 n3736 VSS VSS nmos w=1u l=1u
M7573 n3738 n3742 net2293 VDD pmos w=2u l=1u
M7574 net2293 n3736 VDD VDD pmos w=2u l=1u
M7575 n3742 n2275 VSS VSS nmos w=1u l=1u
M7576 n3742 n3743 VSS VSS nmos w=1u l=1u
M7577 n3742 n2275 net2294 VDD pmos w=2u l=1u
M7578 net2294 n3743 VDD VDD pmos w=2u l=1u
M7579 n2275 N256 VDD VDD pmos w=2u l=1u
M7580 n2275 N256 VSS VSS nmos w=1u l=1u
M7581 n3743 n3745 VSS VSS nmos w=1u l=1u
M7582 n3743 n3744 VSS VSS nmos w=1u l=1u
M7583 n3743 n3745 net2295 VDD pmos w=2u l=1u
M7584 net2295 n3744 VDD VDD pmos w=2u l=1u
M7585 n3744 n3746 VSS VSS nmos w=1u l=1u
M7586 n3744 N239 VSS VSS nmos w=1u l=1u
M7587 n3744 n3746 net2296 VDD pmos w=2u l=1u
M7588 net2296 N239 VDD VDD pmos w=2u l=1u
M7589 n3730 net2297 VSS VSS nmos w=1u l=1u
M7590 net2298 n3748 VSS VSS nmos w=1u l=1u
M7591 net2297 n3747 net2298 VSS nmos w=1u l=1u
M7592 net2297 n3748 VDD VDD pmos w=2u l=1u
M7593 net2297 n3747 VDD VDD pmos w=2u l=1u
M7594 n3730 net2297 VDD VDD pmos w=2u l=1u
M7595 n3723 n3720 VSS VSS nmos w=1u l=1u
M7596 n3723 n3721 VSS VSS nmos w=1u l=1u
M7597 n3723 n3720 net2299 VDD pmos w=2u l=1u
M7598 net2299 n3721 VDD VDD pmos w=2u l=1u
M7599 n3720 n3749 VDD VDD pmos w=2u l=1u
M7600 n3720 n3749 VSS VSS nmos w=1u l=1u
M7601 n3715 n3751 VSS VSS nmos w=1u l=1u
M7602 n3715 n3750 VSS VSS nmos w=1u l=1u
M7603 n3715 n3751 net2300 VDD pmos w=2u l=1u
M7604 net2300 n3750 VDD VDD pmos w=2u l=1u
M7605 n3751 net2301 VSS VSS nmos w=1u l=1u
M7606 net2302 n3712 VSS VSS nmos w=1u l=1u
M7607 net2301 n3713 net2302 VSS nmos w=1u l=1u
M7608 net2301 n3712 VDD VDD pmos w=2u l=1u
M7609 net2301 n3713 VDD VDD pmos w=2u l=1u
M7610 n3751 net2301 VDD VDD pmos w=2u l=1u
M7611 n3750 n3711 VDD VDD pmos w=2u l=1u
M7612 n3750 n3711 VSS VSS nmos w=1u l=1u
M7613 n3705 n3753 VSS VSS nmos w=1u l=1u
M7614 n3705 n3752 VSS VSS nmos w=1u l=1u
M7615 n3705 n3753 net2303 VDD pmos w=2u l=1u
M7616 net2303 n3752 VDD VDD pmos w=2u l=1u
M7617 n3753 n3702 VSS VSS nmos w=1u l=1u
M7618 n3753 n3703 VSS VSS nmos w=1u l=1u
M7619 n3753 n3702 net2304 VDD pmos w=2u l=1u
M7620 net2304 n3703 VDD VDD pmos w=2u l=1u
M7621 n3752 n3701 VDD VDD pmos w=2u l=1u
M7622 n3752 n3701 VSS VSS nmos w=1u l=1u
M7623 n3695 n3755 VSS VSS nmos w=1u l=1u
M7624 n3695 n3754 VSS VSS nmos w=1u l=1u
M7625 n3695 n3755 net2305 VDD pmos w=2u l=1u
M7626 net2305 n3754 VDD VDD pmos w=2u l=1u
M7627 n3755 n3692 VSS VSS nmos w=1u l=1u
M7628 n3755 n3693 VSS VSS nmos w=1u l=1u
M7629 n3755 n3692 net2306 VDD pmos w=2u l=1u
M7630 net2306 n3693 VDD VDD pmos w=2u l=1u
M7631 n3754 n3691 VDD VDD pmos w=2u l=1u
M7632 n3754 n3691 VSS VSS nmos w=1u l=1u
M7633 n3685 n3757 VSS VSS nmos w=1u l=1u
M7634 n3685 n3756 VSS VSS nmos w=1u l=1u
M7635 n3685 n3757 net2307 VDD pmos w=2u l=1u
M7636 net2307 n3756 VDD VDD pmos w=2u l=1u
M7637 n3757 n3682 VSS VSS nmos w=1u l=1u
M7638 n3757 n3683 VSS VSS nmos w=1u l=1u
M7639 n3757 n3682 net2308 VDD pmos w=2u l=1u
M7640 net2308 n3683 VDD VDD pmos w=2u l=1u
M7641 n3756 n3681 VDD VDD pmos w=2u l=1u
M7642 n3756 n3681 VSS VSS nmos w=1u l=1u
M7643 n3675 n3759 VSS VSS nmos w=1u l=1u
M7644 n3675 n3758 VSS VSS nmos w=1u l=1u
M7645 n3675 n3759 net2309 VDD pmos w=2u l=1u
M7646 net2309 n3758 VDD VDD pmos w=2u l=1u
M7647 n3759 n3672 VSS VSS nmos w=1u l=1u
M7648 n3759 n3673 VSS VSS nmos w=1u l=1u
M7649 n3759 n3672 net2310 VDD pmos w=2u l=1u
M7650 net2310 n3673 VDD VDD pmos w=2u l=1u
M7651 n3758 n3671 VDD VDD pmos w=2u l=1u
M7652 n3758 n3671 VSS VSS nmos w=1u l=1u
M7653 n3665 n3761 VSS VSS nmos w=1u l=1u
M7654 n3665 n3760 VSS VSS nmos w=1u l=1u
M7655 n3665 n3761 net2311 VDD pmos w=2u l=1u
M7656 net2311 n3760 VDD VDD pmos w=2u l=1u
M7657 n3761 n3662 VSS VSS nmos w=1u l=1u
M7658 n3761 n3663 VSS VSS nmos w=1u l=1u
M7659 n3761 n3662 net2312 VDD pmos w=2u l=1u
M7660 net2312 n3663 VDD VDD pmos w=2u l=1u
M7661 n3760 n3661 VDD VDD pmos w=2u l=1u
M7662 n3760 n3661 VSS VSS nmos w=1u l=1u
M7663 n3655 n3763 VSS VSS nmos w=1u l=1u
M7664 n3655 n3762 VSS VSS nmos w=1u l=1u
M7665 n3655 n3763 net2313 VDD pmos w=2u l=1u
M7666 net2313 n3762 VDD VDD pmos w=2u l=1u
M7667 n3763 n3652 VSS VSS nmos w=1u l=1u
M7668 n3763 n3653 VSS VSS nmos w=1u l=1u
M7669 n3763 n3652 net2314 VDD pmos w=2u l=1u
M7670 net2314 n3653 VDD VDD pmos w=2u l=1u
M7671 n3762 n3651 VDD VDD pmos w=2u l=1u
M7672 n3762 n3651 VSS VSS nmos w=1u l=1u
M7673 n3645 n3765 VSS VSS nmos w=1u l=1u
M7674 n3645 n3764 VSS VSS nmos w=1u l=1u
M7675 n3645 n3765 net2315 VDD pmos w=2u l=1u
M7676 net2315 n3764 VDD VDD pmos w=2u l=1u
M7677 n3765 n3642 VSS VSS nmos w=1u l=1u
M7678 n3765 n3643 VSS VSS nmos w=1u l=1u
M7679 n3765 n3642 net2316 VDD pmos w=2u l=1u
M7680 net2316 n3643 VDD VDD pmos w=2u l=1u
M7681 n3764 n3641 VDD VDD pmos w=2u l=1u
M7682 n3764 n3641 VSS VSS nmos w=1u l=1u
M7683 n3635 n3767 VSS VSS nmos w=1u l=1u
M7684 n3635 n3766 VSS VSS nmos w=1u l=1u
M7685 n3635 n3767 net2317 VDD pmos w=2u l=1u
M7686 net2317 n3766 VDD VDD pmos w=2u l=1u
M7687 n3767 n3632 VSS VSS nmos w=1u l=1u
M7688 n3767 n3633 VSS VSS nmos w=1u l=1u
M7689 n3767 n3632 net2318 VDD pmos w=2u l=1u
M7690 net2318 n3633 VDD VDD pmos w=2u l=1u
M7691 n3766 n3631 VDD VDD pmos w=2u l=1u
M7692 n3766 n3631 VSS VSS nmos w=1u l=1u
M7693 n3624 n3769 VSS VSS nmos w=1u l=1u
M7694 n3624 n3768 VSS VSS nmos w=1u l=1u
M7695 n3624 n3769 net2319 VDD pmos w=2u l=1u
M7696 net2319 n3768 VDD VDD pmos w=2u l=1u
M7697 n3769 n3622 VSS VSS nmos w=1u l=1u
M7698 n3769 n3623 VSS VSS nmos w=1u l=1u
M7699 n3769 n3622 net2320 VDD pmos w=2u l=1u
M7700 net2320 n3623 VDD VDD pmos w=2u l=1u
M7701 n3768 n3621 VDD VDD pmos w=2u l=1u
M7702 n3768 n3621 VSS VSS nmos w=1u l=1u
M7703 n3614 net2321 VSS VSS nmos w=1u l=1u
M7704 net2322 n3612 VSS VSS nmos w=1u l=1u
M7705 net2321 n3613 net2322 VSS nmos w=1u l=1u
M7706 net2321 n3612 VDD VDD pmos w=2u l=1u
M7707 net2321 n3613 VDD VDD pmos w=2u l=1u
M7708 n3614 net2321 VDD VDD pmos w=2u l=1u
M7709 N5971 n3770 net2323 VSS nmos w=1u l=1u
M7710 net2323 n3612 VSS VSS nmos w=1u l=1u
M7711 N5971 n3770 VDD VDD pmos w=2u l=1u
M7712 N5971 n3612 VDD VDD pmos w=2u l=1u
M7713 n3770 N1 net2324 VSS nmos w=1u l=1u
M7714 net2324 n3771 VSS VSS nmos w=1u l=1u
M7715 n3770 N1 VDD VDD pmos w=2u l=1u
M7716 n3770 n3771 VDD VDD pmos w=2u l=1u
M7717 n3771 n2232 VSS VSS nmos w=1u l=1u
M7718 n3771 n3772 VSS VSS nmos w=1u l=1u
M7719 n3771 n2232 net2325 VDD pmos w=2u l=1u
M7720 net2325 n3772 VDD VDD pmos w=2u l=1u
M7721 n2232 N511 VDD VDD pmos w=2u l=1u
M7722 n2232 N511 VSS VSS nmos w=1u l=1u
M7723 n3612 n3773 net2326 VSS nmos w=1u l=1u
M7724 net2326 n3772 VSS VSS nmos w=1u l=1u
M7725 n3612 n3773 VDD VDD pmos w=2u l=1u
M7726 n3612 n3772 VDD VDD pmos w=2u l=1u
M7727 n3773 N511 net2327 VSS nmos w=1u l=1u
M7728 net2327 N1 VSS VSS nmos w=1u l=1u
M7729 n3773 N511 VDD VDD pmos w=2u l=1u
M7730 n3773 N1 VDD VDD pmos w=2u l=1u
M7731 n3772 net2328 VSS VSS nmos w=1u l=1u
M7732 net2329 n3613 VSS VSS nmos w=1u l=1u
M7733 net2328 n3774 net2329 VSS nmos w=1u l=1u
M7734 net2328 n3613 VDD VDD pmos w=2u l=1u
M7735 net2328 n3774 VDD VDD pmos w=2u l=1u
M7736 n3772 net2328 VDD VDD pmos w=2u l=1u
M7737 n3613 n3776 net2330 VSS nmos w=1u l=1u
M7738 net2330 n3775 VSS VSS nmos w=1u l=1u
M7739 n3613 n3776 VDD VDD pmos w=2u l=1u
M7740 n3613 n3775 VDD VDD pmos w=2u l=1u
M7741 n3776 n3778 net2331 VSS nmos w=1u l=1u
M7742 net2331 n3777 VSS VSS nmos w=1u l=1u
M7743 n3776 n3778 VDD VDD pmos w=2u l=1u
M7744 n3776 n3777 VDD VDD pmos w=2u l=1u
M7745 n3777 net2332 VSS VSS nmos w=1u l=1u
M7746 net2332 n3779 VSS VSS nmos w=1u l=1u
M7747 net2332 n3780 VSS VSS nmos w=1u l=1u
M7748 net2332 n3780 net2333 VDD pmos w=2u l=1u
M7749 n3777 net2332 VDD VDD pmos w=2u l=1u
M7750 net2333 n3779 VDD VDD pmos w=2u l=1u
M7751 net2334 n3622 VSS VSS nmos w=1u l=1u
M7752 net2335 n3623 VSS VSS nmos w=1u l=1u
M7753 n3775 net2336 VSS VSS nmos w=1u l=1u
M7754 net2336 n3622 net2337 VSS nmos w=1u l=1u
M7755 net2336 net2334 net2335 VSS nmos w=1u l=1u
M7756 net2337 net2335 VSS VSS nmos w=1u l=1u
M7757 net2336 net2334 net2338 VDD pmos w=2u l=1u
M7758 net2334 n3622 VDD VDD pmos w=2u l=1u
M7759 net2335 n3622 net2336 VDD pmos w=2u l=1u
M7760 net2335 n3623 VDD VDD pmos w=2u l=1u
M7761 n3775 net2336 VDD VDD pmos w=2u l=1u
M7762 net2338 net2335 VDD VDD pmos w=2u l=1u
M7763 n3774 n3782 net2339 VSS nmos w=1u l=1u
M7764 net2339 n3781 VSS VSS nmos w=1u l=1u
M7765 n3774 n3782 VDD VDD pmos w=2u l=1u
M7766 n3774 n3781 VDD VDD pmos w=2u l=1u
M7767 net2340 n3623 VSS VSS nmos w=1u l=1u
M7768 net2341 n3783 VSS VSS nmos w=1u l=1u
M7769 n3782 net2342 VSS VSS nmos w=1u l=1u
M7770 net2342 n3623 net2343 VSS nmos w=1u l=1u
M7771 net2342 net2340 net2341 VSS nmos w=1u l=1u
M7772 net2343 net2341 VSS VSS nmos w=1u l=1u
M7773 net2342 net2340 net2344 VDD pmos w=2u l=1u
M7774 net2340 n3623 VDD VDD pmos w=2u l=1u
M7775 net2341 n3623 net2342 VDD pmos w=2u l=1u
M7776 net2341 n3783 VDD VDD pmos w=2u l=1u
M7777 n3782 net2342 VDD VDD pmos w=2u l=1u
M7778 net2344 net2341 VDD VDD pmos w=2u l=1u
M7779 n3623 n2271 VSS VSS nmos w=1u l=1u
M7780 n3623 n3603 VSS VSS nmos w=1u l=1u
M7781 n3623 n2271 net2345 VDD pmos w=2u l=1u
M7782 net2345 n3603 VDD VDD pmos w=2u l=1u
M7783 n3783 n3622 VDD VDD pmos w=2u l=1u
M7784 n3783 n3622 VSS VSS nmos w=1u l=1u
M7785 n3622 n3621 net2346 VSS nmos w=1u l=1u
M7786 net2346 n3784 VSS VSS nmos w=1u l=1u
M7787 n3622 n3621 VDD VDD pmos w=2u l=1u
M7788 n3622 n3784 VDD VDD pmos w=2u l=1u
M7789 n3621 n3786 net2347 VSS nmos w=1u l=1u
M7790 net2347 n3785 VSS VSS nmos w=1u l=1u
M7791 n3621 n3786 VDD VDD pmos w=2u l=1u
M7792 n3621 n3785 VDD VDD pmos w=2u l=1u
M7793 n3786 n3788 net2348 VSS nmos w=1u l=1u
M7794 net2348 n3787 VSS VSS nmos w=1u l=1u
M7795 n3786 n3788 VDD VDD pmos w=2u l=1u
M7796 n3786 n3787 VDD VDD pmos w=2u l=1u
M7797 n3787 n3790 net2349 VSS nmos w=1u l=1u
M7798 net2349 n3789 VSS VSS nmos w=1u l=1u
M7799 n3787 n3790 VDD VDD pmos w=2u l=1u
M7800 n3787 n3789 VDD VDD pmos w=2u l=1u
M7801 net2350 n3632 VSS VSS nmos w=1u l=1u
M7802 net2351 n3633 VSS VSS nmos w=1u l=1u
M7803 n3785 net2352 VSS VSS nmos w=1u l=1u
M7804 net2352 n3632 net2353 VSS nmos w=1u l=1u
M7805 net2352 net2350 net2351 VSS nmos w=1u l=1u
M7806 net2353 net2351 VSS VSS nmos w=1u l=1u
M7807 net2352 net2350 net2354 VDD pmos w=2u l=1u
M7808 net2350 n3632 VDD VDD pmos w=2u l=1u
M7809 net2351 n3632 net2352 VDD pmos w=2u l=1u
M7810 net2351 n3633 VDD VDD pmos w=2u l=1u
M7811 n3785 net2352 VDD VDD pmos w=2u l=1u
M7812 net2354 net2351 VDD VDD pmos w=2u l=1u
M7813 n3784 n3792 net2355 VSS nmos w=1u l=1u
M7814 net2355 n3791 VSS VSS nmos w=1u l=1u
M7815 n3784 n3792 VDD VDD pmos w=2u l=1u
M7816 n3784 n3791 VDD VDD pmos w=2u l=1u
M7817 net2356 n3633 VSS VSS nmos w=1u l=1u
M7818 net2357 n3793 VSS VSS nmos w=1u l=1u
M7819 n3792 net2358 VSS VSS nmos w=1u l=1u
M7820 net2358 n3633 net2359 VSS nmos w=1u l=1u
M7821 net2358 net2356 net2357 VSS nmos w=1u l=1u
M7822 net2359 net2357 VSS VSS nmos w=1u l=1u
M7823 net2358 net2356 net2360 VDD pmos w=2u l=1u
M7824 net2356 n3633 VDD VDD pmos w=2u l=1u
M7825 net2357 n3633 net2358 VDD pmos w=2u l=1u
M7826 net2357 n3793 VDD VDD pmos w=2u l=1u
M7827 n3792 net2358 VDD VDD pmos w=2u l=1u
M7828 net2360 net2357 VDD VDD pmos w=2u l=1u
M7829 n3633 n2321 VSS VSS nmos w=1u l=1u
M7830 n3633 n3456 VSS VSS nmos w=1u l=1u
M7831 n3633 n2321 net2361 VDD pmos w=2u l=1u
M7832 net2361 n3456 VDD VDD pmos w=2u l=1u
M7833 n3793 n3632 VDD VDD pmos w=2u l=1u
M7834 n3793 n3632 VSS VSS nmos w=1u l=1u
M7835 n3632 n3631 net2362 VSS nmos w=1u l=1u
M7836 net2362 n3794 VSS VSS nmos w=1u l=1u
M7837 n3632 n3631 VDD VDD pmos w=2u l=1u
M7838 n3632 n3794 VDD VDD pmos w=2u l=1u
M7839 n3631 n3796 net2363 VSS nmos w=1u l=1u
M7840 net2363 n3795 VSS VSS nmos w=1u l=1u
M7841 n3631 n3796 VDD VDD pmos w=2u l=1u
M7842 n3631 n3795 VDD VDD pmos w=2u l=1u
M7843 n3796 n3798 net2364 VSS nmos w=1u l=1u
M7844 net2364 n3797 VSS VSS nmos w=1u l=1u
M7845 n3796 n3798 VDD VDD pmos w=2u l=1u
M7846 n3796 n3797 VDD VDD pmos w=2u l=1u
M7847 n3797 n3800 net2365 VSS nmos w=1u l=1u
M7848 net2365 n3799 VSS VSS nmos w=1u l=1u
M7849 n3797 n3800 VDD VDD pmos w=2u l=1u
M7850 n3797 n3799 VDD VDD pmos w=2u l=1u
M7851 net2366 n3642 VSS VSS nmos w=1u l=1u
M7852 net2367 n3643 VSS VSS nmos w=1u l=1u
M7853 n3795 net2368 VSS VSS nmos w=1u l=1u
M7854 net2368 n3642 net2369 VSS nmos w=1u l=1u
M7855 net2368 net2366 net2367 VSS nmos w=1u l=1u
M7856 net2369 net2367 VSS VSS nmos w=1u l=1u
M7857 net2368 net2366 net2370 VDD pmos w=2u l=1u
M7858 net2366 n3642 VDD VDD pmos w=2u l=1u
M7859 net2367 n3642 net2368 VDD pmos w=2u l=1u
M7860 net2367 n3643 VDD VDD pmos w=2u l=1u
M7861 n3795 net2368 VDD VDD pmos w=2u l=1u
M7862 net2370 net2367 VDD VDD pmos w=2u l=1u
M7863 n3643 n3801 VDD VDD pmos w=2u l=1u
M7864 n3643 n3801 VSS VSS nmos w=1u l=1u
M7865 n3794 n3803 net2371 VSS nmos w=1u l=1u
M7866 net2371 n3802 VSS VSS nmos w=1u l=1u
M7867 n3794 n3803 VDD VDD pmos w=2u l=1u
M7868 n3794 n3802 VDD VDD pmos w=2u l=1u
M7869 net2372 n3801 VSS VSS nmos w=1u l=1u
M7870 net2373 n3642 VSS VSS nmos w=1u l=1u
M7871 n3803 net2374 VSS VSS nmos w=1u l=1u
M7872 net2374 n3801 net2375 VSS nmos w=1u l=1u
M7873 net2374 net2372 net2373 VSS nmos w=1u l=1u
M7874 net2375 net2373 VSS VSS nmos w=1u l=1u
M7875 net2374 net2372 net2376 VDD pmos w=2u l=1u
M7876 net2372 n3801 VDD VDD pmos w=2u l=1u
M7877 net2373 n3801 net2374 VDD pmos w=2u l=1u
M7878 net2373 n3642 VDD VDD pmos w=2u l=1u
M7879 n3803 net2374 VDD VDD pmos w=2u l=1u
M7880 net2376 net2373 VDD VDD pmos w=2u l=1u
M7881 n3801 N460 net2377 VSS nmos w=1u l=1u
M7882 net2377 N52 VSS VSS nmos w=1u l=1u
M7883 n3801 N460 VDD VDD pmos w=2u l=1u
M7884 n3801 N52 VDD VDD pmos w=2u l=1u
M7885 n3642 n3641 net2378 VSS nmos w=1u l=1u
M7886 net2378 n3804 VSS VSS nmos w=1u l=1u
M7887 n3642 n3641 VDD VDD pmos w=2u l=1u
M7888 n3642 n3804 VDD VDD pmos w=2u l=1u
M7889 n3641 n3806 net2379 VSS nmos w=1u l=1u
M7890 net2379 n3805 VSS VSS nmos w=1u l=1u
M7891 n3641 n3806 VDD VDD pmos w=2u l=1u
M7892 n3641 n3805 VDD VDD pmos w=2u l=1u
M7893 n3806 n3808 net2380 VSS nmos w=1u l=1u
M7894 net2380 n3807 VSS VSS nmos w=1u l=1u
M7895 n3806 n3808 VDD VDD pmos w=2u l=1u
M7896 n3806 n3807 VDD VDD pmos w=2u l=1u
M7897 n3807 n3810 net2381 VSS nmos w=1u l=1u
M7898 net2381 n3809 VSS VSS nmos w=1u l=1u
M7899 n3807 n3810 VDD VDD pmos w=2u l=1u
M7900 n3807 n3809 VDD VDD pmos w=2u l=1u
M7901 net2382 n3652 VSS VSS nmos w=1u l=1u
M7902 net2383 n3653 VSS VSS nmos w=1u l=1u
M7903 n3805 net2384 VSS VSS nmos w=1u l=1u
M7904 net2384 n3652 net2385 VSS nmos w=1u l=1u
M7905 net2384 net2382 net2383 VSS nmos w=1u l=1u
M7906 net2385 net2383 VSS VSS nmos w=1u l=1u
M7907 net2384 net2382 net2386 VDD pmos w=2u l=1u
M7908 net2382 n3652 VDD VDD pmos w=2u l=1u
M7909 net2383 n3652 net2384 VDD pmos w=2u l=1u
M7910 net2383 n3653 VDD VDD pmos w=2u l=1u
M7911 n3805 net2384 VDD VDD pmos w=2u l=1u
M7912 net2386 net2383 VDD VDD pmos w=2u l=1u
M7913 n3653 n3811 VDD VDD pmos w=2u l=1u
M7914 n3653 n3811 VSS VSS nmos w=1u l=1u
M7915 n3804 n3813 net2387 VSS nmos w=1u l=1u
M7916 net2387 n3812 VSS VSS nmos w=1u l=1u
M7917 n3804 n3813 VDD VDD pmos w=2u l=1u
M7918 n3804 n3812 VDD VDD pmos w=2u l=1u
M7919 net2388 n3811 VSS VSS nmos w=1u l=1u
M7920 net2389 n3652 VSS VSS nmos w=1u l=1u
M7921 n3813 net2390 VSS VSS nmos w=1u l=1u
M7922 net2390 n3811 net2391 VSS nmos w=1u l=1u
M7923 net2390 net2388 net2389 VSS nmos w=1u l=1u
M7924 net2391 net2389 VSS VSS nmos w=1u l=1u
M7925 net2390 net2388 net2392 VDD pmos w=2u l=1u
M7926 net2388 n3811 VDD VDD pmos w=2u l=1u
M7927 net2389 n3811 net2390 VDD pmos w=2u l=1u
M7928 net2389 n3652 VDD VDD pmos w=2u l=1u
M7929 n3813 net2390 VDD VDD pmos w=2u l=1u
M7930 net2392 net2389 VDD VDD pmos w=2u l=1u
M7931 n3811 N443 net2393 VSS nmos w=1u l=1u
M7932 net2393 N69 VSS VSS nmos w=1u l=1u
M7933 n3811 N443 VDD VDD pmos w=2u l=1u
M7934 n3811 N69 VDD VDD pmos w=2u l=1u
M7935 n3652 n3651 net2394 VSS nmos w=1u l=1u
M7936 net2394 n3814 VSS VSS nmos w=1u l=1u
M7937 n3652 n3651 VDD VDD pmos w=2u l=1u
M7938 n3652 n3814 VDD VDD pmos w=2u l=1u
M7939 n3651 n3816 net2395 VSS nmos w=1u l=1u
M7940 net2395 n3815 VSS VSS nmos w=1u l=1u
M7941 n3651 n3816 VDD VDD pmos w=2u l=1u
M7942 n3651 n3815 VDD VDD pmos w=2u l=1u
M7943 n3816 n3818 net2396 VSS nmos w=1u l=1u
M7944 net2396 n3817 VSS VSS nmos w=1u l=1u
M7945 n3816 n3818 VDD VDD pmos w=2u l=1u
M7946 n3816 n3817 VDD VDD pmos w=2u l=1u
M7947 n3817 n3820 net2397 VSS nmos w=1u l=1u
M7948 net2397 n3819 VSS VSS nmos w=1u l=1u
M7949 n3817 n3820 VDD VDD pmos w=2u l=1u
M7950 n3817 n3819 VDD VDD pmos w=2u l=1u
M7951 net2398 n3662 VSS VSS nmos w=1u l=1u
M7952 net2399 n3663 VSS VSS nmos w=1u l=1u
M7953 n3815 net2400 VSS VSS nmos w=1u l=1u
M7954 net2400 n3662 net2401 VSS nmos w=1u l=1u
M7955 net2400 net2398 net2399 VSS nmos w=1u l=1u
M7956 net2401 net2399 VSS VSS nmos w=1u l=1u
M7957 net2400 net2398 net2402 VDD pmos w=2u l=1u
M7958 net2398 n3662 VDD VDD pmos w=2u l=1u
M7959 net2399 n3662 net2400 VDD pmos w=2u l=1u
M7960 net2399 n3663 VDD VDD pmos w=2u l=1u
M7961 n3815 net2400 VDD VDD pmos w=2u l=1u
M7962 net2402 net2399 VDD VDD pmos w=2u l=1u
M7963 n3663 n3821 VDD VDD pmos w=2u l=1u
M7964 n3663 n3821 VSS VSS nmos w=1u l=1u
M7965 n3814 n3823 net2403 VSS nmos w=1u l=1u
M7966 net2403 n3822 VSS VSS nmos w=1u l=1u
M7967 n3814 n3823 VDD VDD pmos w=2u l=1u
M7968 n3814 n3822 VDD VDD pmos w=2u l=1u
M7969 net2404 n3821 VSS VSS nmos w=1u l=1u
M7970 net2405 n3662 VSS VSS nmos w=1u l=1u
M7971 n3823 net2406 VSS VSS nmos w=1u l=1u
M7972 net2406 n3821 net2407 VSS nmos w=1u l=1u
M7973 net2406 net2404 net2405 VSS nmos w=1u l=1u
M7974 net2407 net2405 VSS VSS nmos w=1u l=1u
M7975 net2406 net2404 net2408 VDD pmos w=2u l=1u
M7976 net2404 n3821 VDD VDD pmos w=2u l=1u
M7977 net2405 n3821 net2406 VDD pmos w=2u l=1u
M7978 net2405 n3662 VDD VDD pmos w=2u l=1u
M7979 n3823 net2406 VDD VDD pmos w=2u l=1u
M7980 net2408 net2405 VDD VDD pmos w=2u l=1u
M7981 n3821 N426 net2409 VSS nmos w=1u l=1u
M7982 net2409 N86 VSS VSS nmos w=1u l=1u
M7983 n3821 N426 VDD VDD pmos w=2u l=1u
M7984 n3821 N86 VDD VDD pmos w=2u l=1u
M7985 n3662 n3661 net2410 VSS nmos w=1u l=1u
M7986 net2410 n3824 VSS VSS nmos w=1u l=1u
M7987 n3662 n3661 VDD VDD pmos w=2u l=1u
M7988 n3662 n3824 VDD VDD pmos w=2u l=1u
M7989 n3661 n3826 net2411 VSS nmos w=1u l=1u
M7990 net2411 n3825 VSS VSS nmos w=1u l=1u
M7991 n3661 n3826 VDD VDD pmos w=2u l=1u
M7992 n3661 n3825 VDD VDD pmos w=2u l=1u
M7993 n3826 n3828 net2412 VSS nmos w=1u l=1u
M7994 net2412 n3827 VSS VSS nmos w=1u l=1u
M7995 n3826 n3828 VDD VDD pmos w=2u l=1u
M7996 n3826 n3827 VDD VDD pmos w=2u l=1u
M7997 n3827 n3830 net2413 VSS nmos w=1u l=1u
M7998 net2413 n3829 VSS VSS nmos w=1u l=1u
M7999 n3827 n3830 VDD VDD pmos w=2u l=1u
M8000 n3827 n3829 VDD VDD pmos w=2u l=1u
M8001 net2414 n3672 VSS VSS nmos w=1u l=1u
M8002 net2415 n3673 VSS VSS nmos w=1u l=1u
M8003 n3825 net2416 VSS VSS nmos w=1u l=1u
M8004 net2416 n3672 net2417 VSS nmos w=1u l=1u
M8005 net2416 net2414 net2415 VSS nmos w=1u l=1u
M8006 net2417 net2415 VSS VSS nmos w=1u l=1u
M8007 net2416 net2414 net2418 VDD pmos w=2u l=1u
M8008 net2414 n3672 VDD VDD pmos w=2u l=1u
M8009 net2415 n3672 net2416 VDD pmos w=2u l=1u
M8010 net2415 n3673 VDD VDD pmos w=2u l=1u
M8011 n3825 net2416 VDD VDD pmos w=2u l=1u
M8012 net2418 net2415 VDD VDD pmos w=2u l=1u
M8013 n3673 n3831 VDD VDD pmos w=2u l=1u
M8014 n3673 n3831 VSS VSS nmos w=1u l=1u
M8015 n3824 n3833 net2419 VSS nmos w=1u l=1u
M8016 net2419 n3832 VSS VSS nmos w=1u l=1u
M8017 n3824 n3833 VDD VDD pmos w=2u l=1u
M8018 n3824 n3832 VDD VDD pmos w=2u l=1u
M8019 net2420 n3831 VSS VSS nmos w=1u l=1u
M8020 net2421 n3672 VSS VSS nmos w=1u l=1u
M8021 n3833 net2422 VSS VSS nmos w=1u l=1u
M8022 net2422 n3831 net2423 VSS nmos w=1u l=1u
M8023 net2422 net2420 net2421 VSS nmos w=1u l=1u
M8024 net2423 net2421 VSS VSS nmos w=1u l=1u
M8025 net2422 net2420 net2424 VDD pmos w=2u l=1u
M8026 net2420 n3831 VDD VDD pmos w=2u l=1u
M8027 net2421 n3831 net2422 VDD pmos w=2u l=1u
M8028 net2421 n3672 VDD VDD pmos w=2u l=1u
M8029 n3833 net2422 VDD VDD pmos w=2u l=1u
M8030 net2424 net2421 VDD VDD pmos w=2u l=1u
M8031 n3831 N409 net2425 VSS nmos w=1u l=1u
M8032 net2425 N103 VSS VSS nmos w=1u l=1u
M8033 n3831 N409 VDD VDD pmos w=2u l=1u
M8034 n3831 N103 VDD VDD pmos w=2u l=1u
M8035 n3672 n3671 net2426 VSS nmos w=1u l=1u
M8036 net2426 n3834 VSS VSS nmos w=1u l=1u
M8037 n3672 n3671 VDD VDD pmos w=2u l=1u
M8038 n3672 n3834 VDD VDD pmos w=2u l=1u
M8039 n3671 n3836 net2427 VSS nmos w=1u l=1u
M8040 net2427 n3835 VSS VSS nmos w=1u l=1u
M8041 n3671 n3836 VDD VDD pmos w=2u l=1u
M8042 n3671 n3835 VDD VDD pmos w=2u l=1u
M8043 n3836 n3838 net2428 VSS nmos w=1u l=1u
M8044 net2428 n3837 VSS VSS nmos w=1u l=1u
M8045 n3836 n3838 VDD VDD pmos w=2u l=1u
M8046 n3836 n3837 VDD VDD pmos w=2u l=1u
M8047 n3837 n3840 net2429 VSS nmos w=1u l=1u
M8048 net2429 n3839 VSS VSS nmos w=1u l=1u
M8049 n3837 n3840 VDD VDD pmos w=2u l=1u
M8050 n3837 n3839 VDD VDD pmos w=2u l=1u
M8051 net2430 n3682 VSS VSS nmos w=1u l=1u
M8052 net2431 n3683 VSS VSS nmos w=1u l=1u
M8053 n3835 net2432 VSS VSS nmos w=1u l=1u
M8054 net2432 n3682 net2433 VSS nmos w=1u l=1u
M8055 net2432 net2430 net2431 VSS nmos w=1u l=1u
M8056 net2433 net2431 VSS VSS nmos w=1u l=1u
M8057 net2432 net2430 net2434 VDD pmos w=2u l=1u
M8058 net2430 n3682 VDD VDD pmos w=2u l=1u
M8059 net2431 n3682 net2432 VDD pmos w=2u l=1u
M8060 net2431 n3683 VDD VDD pmos w=2u l=1u
M8061 n3835 net2432 VDD VDD pmos w=2u l=1u
M8062 net2434 net2431 VDD VDD pmos w=2u l=1u
M8063 n3683 n3841 VDD VDD pmos w=2u l=1u
M8064 n3683 n3841 VSS VSS nmos w=1u l=1u
M8065 n3834 n3843 net2435 VSS nmos w=1u l=1u
M8066 net2435 n3842 VSS VSS nmos w=1u l=1u
M8067 n3834 n3843 VDD VDD pmos w=2u l=1u
M8068 n3834 n3842 VDD VDD pmos w=2u l=1u
M8069 net2436 n3841 VSS VSS nmos w=1u l=1u
M8070 net2437 n3682 VSS VSS nmos w=1u l=1u
M8071 n3843 net2438 VSS VSS nmos w=1u l=1u
M8072 net2438 n3841 net2439 VSS nmos w=1u l=1u
M8073 net2438 net2436 net2437 VSS nmos w=1u l=1u
M8074 net2439 net2437 VSS VSS nmos w=1u l=1u
M8075 net2438 net2436 net2440 VDD pmos w=2u l=1u
M8076 net2436 n3841 VDD VDD pmos w=2u l=1u
M8077 net2437 n3841 net2438 VDD pmos w=2u l=1u
M8078 net2437 n3682 VDD VDD pmos w=2u l=1u
M8079 n3843 net2438 VDD VDD pmos w=2u l=1u
M8080 net2440 net2437 VDD VDD pmos w=2u l=1u
M8081 n3841 N392 net2441 VSS nmos w=1u l=1u
M8082 net2441 N120 VSS VSS nmos w=1u l=1u
M8083 n3841 N392 VDD VDD pmos w=2u l=1u
M8084 n3841 N120 VDD VDD pmos w=2u l=1u
M8085 n3682 n3681 net2442 VSS nmos w=1u l=1u
M8086 net2442 n3844 VSS VSS nmos w=1u l=1u
M8087 n3682 n3681 VDD VDD pmos w=2u l=1u
M8088 n3682 n3844 VDD VDD pmos w=2u l=1u
M8089 n3681 n3846 net2443 VSS nmos w=1u l=1u
M8090 net2443 n3845 VSS VSS nmos w=1u l=1u
M8091 n3681 n3846 VDD VDD pmos w=2u l=1u
M8092 n3681 n3845 VDD VDD pmos w=2u l=1u
M8093 n3846 n3848 net2444 VSS nmos w=1u l=1u
M8094 net2444 n3847 VSS VSS nmos w=1u l=1u
M8095 n3846 n3848 VDD VDD pmos w=2u l=1u
M8096 n3846 n3847 VDD VDD pmos w=2u l=1u
M8097 n3847 n3850 net2445 VSS nmos w=1u l=1u
M8098 net2445 n3849 VSS VSS nmos w=1u l=1u
M8099 n3847 n3850 VDD VDD pmos w=2u l=1u
M8100 n3847 n3849 VDD VDD pmos w=2u l=1u
M8101 net2446 n3692 VSS VSS nmos w=1u l=1u
M8102 net2447 n3693 VSS VSS nmos w=1u l=1u
M8103 n3845 net2448 VSS VSS nmos w=1u l=1u
M8104 net2448 n3692 net2449 VSS nmos w=1u l=1u
M8105 net2448 net2446 net2447 VSS nmos w=1u l=1u
M8106 net2449 net2447 VSS VSS nmos w=1u l=1u
M8107 net2448 net2446 net2450 VDD pmos w=2u l=1u
M8108 net2446 n3692 VDD VDD pmos w=2u l=1u
M8109 net2447 n3692 net2448 VDD pmos w=2u l=1u
M8110 net2447 n3693 VDD VDD pmos w=2u l=1u
M8111 n3845 net2448 VDD VDD pmos w=2u l=1u
M8112 net2450 net2447 VDD VDD pmos w=2u l=1u
M8113 n3693 n3851 VDD VDD pmos w=2u l=1u
M8114 n3693 n3851 VSS VSS nmos w=1u l=1u
M8115 n3844 n3853 net2451 VSS nmos w=1u l=1u
M8116 net2451 n3852 VSS VSS nmos w=1u l=1u
M8117 n3844 n3853 VDD VDD pmos w=2u l=1u
M8118 n3844 n3852 VDD VDD pmos w=2u l=1u
M8119 net2452 n3851 VSS VSS nmos w=1u l=1u
M8120 net2453 n3692 VSS VSS nmos w=1u l=1u
M8121 n3853 net2454 VSS VSS nmos w=1u l=1u
M8122 net2454 n3851 net2455 VSS nmos w=1u l=1u
M8123 net2454 net2452 net2453 VSS nmos w=1u l=1u
M8124 net2455 net2453 VSS VSS nmos w=1u l=1u
M8125 net2454 net2452 net2456 VDD pmos w=2u l=1u
M8126 net2452 n3851 VDD VDD pmos w=2u l=1u
M8127 net2453 n3851 net2454 VDD pmos w=2u l=1u
M8128 net2453 n3692 VDD VDD pmos w=2u l=1u
M8129 n3853 net2454 VDD VDD pmos w=2u l=1u
M8130 net2456 net2453 VDD VDD pmos w=2u l=1u
M8131 n3851 N375 net2457 VSS nmos w=1u l=1u
M8132 net2457 N137 VSS VSS nmos w=1u l=1u
M8133 n3851 N375 VDD VDD pmos w=2u l=1u
M8134 n3851 N137 VDD VDD pmos w=2u l=1u
M8135 n3692 n3691 net2458 VSS nmos w=1u l=1u
M8136 net2458 n3854 VSS VSS nmos w=1u l=1u
M8137 n3692 n3691 VDD VDD pmos w=2u l=1u
M8138 n3692 n3854 VDD VDD pmos w=2u l=1u
M8139 n3691 n3856 net2459 VSS nmos w=1u l=1u
M8140 net2459 n3855 VSS VSS nmos w=1u l=1u
M8141 n3691 n3856 VDD VDD pmos w=2u l=1u
M8142 n3691 n3855 VDD VDD pmos w=2u l=1u
M8143 n3856 n3858 net2460 VSS nmos w=1u l=1u
M8144 net2460 n3857 VSS VSS nmos w=1u l=1u
M8145 n3856 n3858 VDD VDD pmos w=2u l=1u
M8146 n3856 n3857 VDD VDD pmos w=2u l=1u
M8147 n3857 net2461 VSS VSS nmos w=1u l=1u
M8148 net2461 n3859 VSS VSS nmos w=1u l=1u
M8149 net2461 n3860 VSS VSS nmos w=1u l=1u
M8150 net2461 n3860 net2462 VDD pmos w=2u l=1u
M8151 n3857 net2461 VDD VDD pmos w=2u l=1u
M8152 net2462 n3859 VDD VDD pmos w=2u l=1u
M8153 net2463 n3702 VSS VSS nmos w=1u l=1u
M8154 net2464 n3703 VSS VSS nmos w=1u l=1u
M8155 n3855 net2465 VSS VSS nmos w=1u l=1u
M8156 net2465 n3702 net2466 VSS nmos w=1u l=1u
M8157 net2465 net2463 net2464 VSS nmos w=1u l=1u
M8158 net2466 net2464 VSS VSS nmos w=1u l=1u
M8159 net2465 net2463 net2467 VDD pmos w=2u l=1u
M8160 net2463 n3702 VDD VDD pmos w=2u l=1u
M8161 net2464 n3702 net2465 VDD pmos w=2u l=1u
M8162 net2464 n3703 VDD VDD pmos w=2u l=1u
M8163 n3855 net2465 VDD VDD pmos w=2u l=1u
M8164 net2467 net2464 VDD VDD pmos w=2u l=1u
M8165 n3703 n3861 VDD VDD pmos w=2u l=1u
M8166 n3703 n3861 VSS VSS nmos w=1u l=1u
M8167 n3854 n3863 net2468 VSS nmos w=1u l=1u
M8168 net2468 n3862 VSS VSS nmos w=1u l=1u
M8169 n3854 n3863 VDD VDD pmos w=2u l=1u
M8170 n3854 n3862 VDD VDD pmos w=2u l=1u
M8171 net2469 n3861 VSS VSS nmos w=1u l=1u
M8172 net2470 n3702 VSS VSS nmos w=1u l=1u
M8173 n3863 net2471 VSS VSS nmos w=1u l=1u
M8174 net2471 n3861 net2472 VSS nmos w=1u l=1u
M8175 net2471 net2469 net2470 VSS nmos w=1u l=1u
M8176 net2472 net2470 VSS VSS nmos w=1u l=1u
M8177 net2471 net2469 net2473 VDD pmos w=2u l=1u
M8178 net2469 n3861 VDD VDD pmos w=2u l=1u
M8179 net2470 n3861 net2471 VDD pmos w=2u l=1u
M8180 net2470 n3702 VDD VDD pmos w=2u l=1u
M8181 n3863 net2471 VDD VDD pmos w=2u l=1u
M8182 net2473 net2470 VDD VDD pmos w=2u l=1u
M8183 n3861 N358 net2474 VSS nmos w=1u l=1u
M8184 net2474 N154 VSS VSS nmos w=1u l=1u
M8185 n3861 N358 VDD VDD pmos w=2u l=1u
M8186 n3861 N154 VDD VDD pmos w=2u l=1u
M8187 n3702 n3701 net2475 VSS nmos w=1u l=1u
M8188 net2475 n3864 VSS VSS nmos w=1u l=1u
M8189 n3702 n3701 VDD VDD pmos w=2u l=1u
M8190 n3702 n3864 VDD VDD pmos w=2u l=1u
M8191 n3701 n3866 net2476 VSS nmos w=1u l=1u
M8192 net2476 n3865 VSS VSS nmos w=1u l=1u
M8193 n3701 n3866 VDD VDD pmos w=2u l=1u
M8194 n3701 n3865 VDD VDD pmos w=2u l=1u
M8195 n3866 n3868 net2477 VSS nmos w=1u l=1u
M8196 net2477 n3867 VSS VSS nmos w=1u l=1u
M8197 n3866 n3868 VDD VDD pmos w=2u l=1u
M8198 n3866 n3867 VDD VDD pmos w=2u l=1u
M8199 n3867 n3870 net2478 VSS nmos w=1u l=1u
M8200 net2478 n3869 VSS VSS nmos w=1u l=1u
M8201 n3867 n3870 VDD VDD pmos w=2u l=1u
M8202 n3867 n3869 VDD VDD pmos w=2u l=1u
M8203 net2479 n3712 VSS VSS nmos w=1u l=1u
M8204 net2480 n3713 VSS VSS nmos w=1u l=1u
M8205 n3865 net2481 VSS VSS nmos w=1u l=1u
M8206 net2481 n3712 net2482 VSS nmos w=1u l=1u
M8207 net2481 net2479 net2480 VSS nmos w=1u l=1u
M8208 net2482 net2480 VSS VSS nmos w=1u l=1u
M8209 net2481 net2479 net2483 VDD pmos w=2u l=1u
M8210 net2479 n3712 VDD VDD pmos w=2u l=1u
M8211 net2480 n3712 net2481 VDD pmos w=2u l=1u
M8212 net2480 n3713 VDD VDD pmos w=2u l=1u
M8213 n3865 net2481 VDD VDD pmos w=2u l=1u
M8214 net2483 net2480 VDD VDD pmos w=2u l=1u
M8215 n3712 n3871 VDD VDD pmos w=2u l=1u
M8216 n3712 n3871 VSS VSS nmos w=1u l=1u
M8217 n3864 n3873 net2484 VSS nmos w=1u l=1u
M8218 net2484 n3872 VSS VSS nmos w=1u l=1u
M8219 n3864 n3873 VDD VDD pmos w=2u l=1u
M8220 n3864 n3872 VDD VDD pmos w=2u l=1u
M8221 net2485 n3713 VSS VSS nmos w=1u l=1u
M8222 net2486 n3871 VSS VSS nmos w=1u l=1u
M8223 n3873 net2487 VSS VSS nmos w=1u l=1u
M8224 net2487 n3713 net2488 VSS nmos w=1u l=1u
M8225 net2487 net2485 net2486 VSS nmos w=1u l=1u
M8226 net2488 net2486 VSS VSS nmos w=1u l=1u
M8227 net2487 net2485 net2489 VDD pmos w=2u l=1u
M8228 net2485 n3713 VDD VDD pmos w=2u l=1u
M8229 net2486 n3713 net2487 VDD pmos w=2u l=1u
M8230 net2486 n3871 VDD VDD pmos w=2u l=1u
M8231 n3873 net2487 VDD VDD pmos w=2u l=1u
M8232 net2489 net2486 VDD VDD pmos w=2u l=1u
M8233 n3713 N341 net2490 VSS nmos w=1u l=1u
M8234 net2490 N171 VSS VSS nmos w=1u l=1u
M8235 n3713 N341 VDD VDD pmos w=2u l=1u
M8236 n3713 N171 VDD VDD pmos w=2u l=1u
M8237 n3871 n3711 net2491 VSS nmos w=1u l=1u
M8238 net2491 n3874 VSS VSS nmos w=1u l=1u
M8239 n3871 n3711 VDD VDD pmos w=2u l=1u
M8240 n3871 n3874 VDD VDD pmos w=2u l=1u
M8241 n3711 n3876 net2492 VSS nmos w=1u l=1u
M8242 net2492 n3875 VSS VSS nmos w=1u l=1u
M8243 n3711 n3876 VDD VDD pmos w=2u l=1u
M8244 n3711 n3875 VDD VDD pmos w=2u l=1u
M8245 n3876 net2493 VSS VSS nmos w=1u l=1u
M8246 net2493 n3877 VSS VSS nmos w=1u l=1u
M8247 net2493 n3878 VSS VSS nmos w=1u l=1u
M8248 net2493 n3878 net2494 VDD pmos w=2u l=1u
M8249 n3876 net2493 VDD VDD pmos w=2u l=1u
M8250 net2494 n3877 VDD VDD pmos w=2u l=1u
M8251 n3875 net2495 VSS VSS nmos w=1u l=1u
M8252 net2496 n3879 VSS VSS nmos w=1u l=1u
M8253 net2495 n3749 net2496 VSS nmos w=1u l=1u
M8254 net2495 n3879 VDD VDD pmos w=2u l=1u
M8255 net2495 n3749 VDD VDD pmos w=2u l=1u
M8256 n3875 net2495 VDD VDD pmos w=2u l=1u
M8257 n3874 n3881 net2497 VSS nmos w=1u l=1u
M8258 net2497 n3880 VSS VSS nmos w=1u l=1u
M8259 n3874 n3881 VDD VDD pmos w=2u l=1u
M8260 n3874 n3880 VDD VDD pmos w=2u l=1u
M8261 n3881 n3749 net2498 VSS nmos w=1u l=1u
M8262 net2498 n3879 VSS VSS nmos w=1u l=1u
M8263 n3881 n3749 VDD VDD pmos w=2u l=1u
M8264 n3881 n3879 VDD VDD pmos w=2u l=1u
M8265 n3749 n3883 net2499 VSS nmos w=1u l=1u
M8266 net2499 n3882 VSS VSS nmos w=1u l=1u
M8267 n3749 n3883 VDD VDD pmos w=2u l=1u
M8268 n3749 n3882 VDD VDD pmos w=2u l=1u
M8269 n3883 N324 net2500 VSS nmos w=1u l=1u
M8270 net2500 N188 VSS VSS nmos w=1u l=1u
M8271 n3883 N324 VDD VDD pmos w=2u l=1u
M8272 n3883 N188 VDD VDD pmos w=2u l=1u
M8273 n3879 N188 net2501 VSS nmos w=1u l=1u
M8274 net2501 n3884 VSS VSS nmos w=1u l=1u
M8275 n3879 N188 VDD VDD pmos w=2u l=1u
M8276 n3879 n3884 VDD VDD pmos w=2u l=1u
M8277 n3884 n3257 VSS VSS nmos w=1u l=1u
M8278 n3884 n3882 VSS VSS nmos w=1u l=1u
M8279 n3884 n3257 net2502 VDD pmos w=2u l=1u
M8280 net2502 n3882 VDD VDD pmos w=2u l=1u
M8281 n3882 n3721 VSS VSS nmos w=1u l=1u
M8282 n3882 n3885 VSS VSS nmos w=1u l=1u
M8283 n3882 n3721 net2503 VDD pmos w=2u l=1u
M8284 net2503 n3885 VDD VDD pmos w=2u l=1u
M8285 n3721 n3887 VSS VSS nmos w=1u l=1u
M8286 n3721 n3886 VSS VSS nmos w=1u l=1u
M8287 n3721 n3887 net2504 VDD pmos w=2u l=1u
M8288 net2504 n3886 VDD VDD pmos w=2u l=1u
M8289 n3885 net2505 VSS VSS nmos w=1u l=1u
M8290 net2506 n3886 VSS VSS nmos w=1u l=1u
M8291 net2505 n3887 net2506 VSS nmos w=1u l=1u
M8292 net2505 n3886 VDD VDD pmos w=2u l=1u
M8293 net2505 n3887 VDD VDD pmos w=2u l=1u
M8294 n3885 net2505 VDD VDD pmos w=2u l=1u
M8295 n3886 n3888 net2507 VSS nmos w=1u l=1u
M8296 net2507 n3747 VSS VSS nmos w=1u l=1u
M8297 n3886 n3888 VDD VDD pmos w=2u l=1u
M8298 n3886 n3747 VDD VDD pmos w=2u l=1u
M8299 n3888 N205 net2508 VSS nmos w=1u l=1u
M8300 net2508 n3889 VSS VSS nmos w=1u l=1u
M8301 n3888 N205 VDD VDD pmos w=2u l=1u
M8302 n3888 n3889 VDD VDD pmos w=2u l=1u
M8303 n3889 n3411 VSS VSS nmos w=1u l=1u
M8304 n3889 n3890 VSS VSS nmos w=1u l=1u
M8305 n3889 n3411 net2509 VDD pmos w=2u l=1u
M8306 net2509 n3890 VDD VDD pmos w=2u l=1u
M8307 n3747 n3891 net2510 VSS nmos w=1u l=1u
M8308 net2510 n3890 VSS VSS nmos w=1u l=1u
M8309 n3747 n3891 VDD VDD pmos w=2u l=1u
M8310 n3747 n3890 VDD VDD pmos w=2u l=1u
M8311 n3891 N307 net2511 VSS nmos w=1u l=1u
M8312 net2511 N205 VSS VSS nmos w=1u l=1u
M8313 n3891 N307 VDD VDD pmos w=2u l=1u
M8314 n3891 N205 VDD VDD pmos w=2u l=1u
M8315 n3890 net2512 VSS VSS nmos w=1u l=1u
M8316 net2513 n3892 VSS VSS nmos w=1u l=1u
M8317 net2512 n3748 net2513 VSS nmos w=1u l=1u
M8318 net2512 n3892 VDD VDD pmos w=2u l=1u
M8319 net2512 n3748 VDD VDD pmos w=2u l=1u
M8320 n3890 net2512 VDD VDD pmos w=2u l=1u
M8321 n3892 net2514 VSS VSS nmos w=1u l=1u
M8322 net2514 n3893 VSS VSS nmos w=1u l=1u
M8323 net2514 n3736 VSS VSS nmos w=1u l=1u
M8324 net2514 n3736 net2515 VDD pmos w=2u l=1u
M8325 n3892 net2514 VDD VDD pmos w=2u l=1u
M8326 net2515 n3893 VDD VDD pmos w=2u l=1u
M8327 n3736 n3894 VDD VDD pmos w=2u l=1u
M8328 n3736 n3894 VSS VSS nmos w=1u l=1u
M8329 n3748 n3895 net2516 VSS nmos w=1u l=1u
M8330 net2516 n3893 VSS VSS nmos w=1u l=1u
M8331 n3748 n3895 VDD VDD pmos w=2u l=1u
M8332 n3748 n3893 VDD VDD pmos w=2u l=1u
M8333 n3895 n3894 net2517 VSS nmos w=1u l=1u
M8334 net2517 n3896 VSS VSS nmos w=1u l=1u
M8335 n3895 n3894 VDD VDD pmos w=2u l=1u
M8336 n3895 n3896 VDD VDD pmos w=2u l=1u
M8337 n3894 N222 net2518 VSS nmos w=1u l=1u
M8338 net2518 n3897 VSS VSS nmos w=1u l=1u
M8339 n3894 N222 VDD VDD pmos w=2u l=1u
M8340 n3894 n3897 VDD VDD pmos w=2u l=1u
M8341 n3897 n3898 VSS VSS nmos w=1u l=1u
M8342 n3897 n2228 VSS VSS nmos w=1u l=1u
M8343 n3897 n3898 net2519 VDD pmos w=2u l=1u
M8344 net2519 n2228 VDD VDD pmos w=2u l=1u
M8345 n2228 N239 VDD VDD pmos w=2u l=1u
M8346 n2228 N239 VSS VSS nmos w=1u l=1u
M8347 n3896 n3900 net2520 VSS nmos w=1u l=1u
M8348 net2520 n3899 VSS VSS nmos w=1u l=1u
M8349 n3896 n3900 VDD VDD pmos w=2u l=1u
M8350 n3896 n3899 VDD VDD pmos w=2u l=1u
M8351 n3900 N239 net2521 VSS nmos w=1u l=1u
M8352 net2521 N273 VSS VSS nmos w=1u l=1u
M8353 n3900 N239 VDD VDD pmos w=2u l=1u
M8354 n3900 N273 VDD VDD pmos w=2u l=1u
M8355 n3899 N290 net2522 VSS nmos w=1u l=1u
M8356 net2522 N222 VSS VSS nmos w=1u l=1u
M8357 n3899 N290 VDD VDD pmos w=2u l=1u
M8358 n3899 N222 VDD VDD pmos w=2u l=1u
M8359 n3887 net2523 VSS VSS nmos w=1u l=1u
M8360 net2524 n3902 VSS VSS nmos w=1u l=1u
M8361 net2523 n3901 net2524 VSS nmos w=1u l=1u
M8362 net2523 n3902 VDD VDD pmos w=2u l=1u
M8363 net2523 n3901 VDD VDD pmos w=2u l=1u
M8364 n3887 net2523 VDD VDD pmos w=2u l=1u
M8365 n3880 n3877 VSS VSS nmos w=1u l=1u
M8366 n3880 n3878 VSS VSS nmos w=1u l=1u
M8367 n3880 n3877 net2525 VDD pmos w=2u l=1u
M8368 net2525 n3878 VDD VDD pmos w=2u l=1u
M8369 n3877 n3903 VDD VDD pmos w=2u l=1u
M8370 n3877 n3903 VSS VSS nmos w=1u l=1u
M8371 n3872 n3905 VSS VSS nmos w=1u l=1u
M8372 n3872 n3904 VSS VSS nmos w=1u l=1u
M8373 n3872 n3905 net2526 VDD pmos w=2u l=1u
M8374 net2526 n3904 VDD VDD pmos w=2u l=1u
M8375 n3905 net2527 VSS VSS nmos w=1u l=1u
M8376 net2528 n3869 VSS VSS nmos w=1u l=1u
M8377 net2527 n3870 net2528 VSS nmos w=1u l=1u
M8378 net2527 n3869 VDD VDD pmos w=2u l=1u
M8379 net2527 n3870 VDD VDD pmos w=2u l=1u
M8380 n3905 net2527 VDD VDD pmos w=2u l=1u
M8381 n3904 n3868 VDD VDD pmos w=2u l=1u
M8382 n3904 n3868 VSS VSS nmos w=1u l=1u
M8383 n3862 n3907 VSS VSS nmos w=1u l=1u
M8384 n3862 n3906 VSS VSS nmos w=1u l=1u
M8385 n3862 n3907 net2529 VDD pmos w=2u l=1u
M8386 net2529 n3906 VDD VDD pmos w=2u l=1u
M8387 n3907 n3859 VSS VSS nmos w=1u l=1u
M8388 n3907 n3860 VSS VSS nmos w=1u l=1u
M8389 n3907 n3859 net2530 VDD pmos w=2u l=1u
M8390 net2530 n3860 VDD VDD pmos w=2u l=1u
M8391 n3906 n3858 VDD VDD pmos w=2u l=1u
M8392 n3906 n3858 VSS VSS nmos w=1u l=1u
M8393 n3852 n3909 VSS VSS nmos w=1u l=1u
M8394 n3852 n3908 VSS VSS nmos w=1u l=1u
M8395 n3852 n3909 net2531 VDD pmos w=2u l=1u
M8396 net2531 n3908 VDD VDD pmos w=2u l=1u
M8397 n3909 net2532 VSS VSS nmos w=1u l=1u
M8398 net2533 n3849 VSS VSS nmos w=1u l=1u
M8399 net2532 n3850 net2533 VSS nmos w=1u l=1u
M8400 net2532 n3849 VDD VDD pmos w=2u l=1u
M8401 net2532 n3850 VDD VDD pmos w=2u l=1u
M8402 n3909 net2532 VDD VDD pmos w=2u l=1u
M8403 n3908 n3848 VDD VDD pmos w=2u l=1u
M8404 n3908 n3848 VSS VSS nmos w=1u l=1u
M8405 n3842 n3911 VSS VSS nmos w=1u l=1u
M8406 n3842 n3910 VSS VSS nmos w=1u l=1u
M8407 n3842 n3911 net2534 VDD pmos w=2u l=1u
M8408 net2534 n3910 VDD VDD pmos w=2u l=1u
M8409 n3911 net2535 VSS VSS nmos w=1u l=1u
M8410 net2536 n3839 VSS VSS nmos w=1u l=1u
M8411 net2535 n3840 net2536 VSS nmos w=1u l=1u
M8412 net2535 n3839 VDD VDD pmos w=2u l=1u
M8413 net2535 n3840 VDD VDD pmos w=2u l=1u
M8414 n3911 net2535 VDD VDD pmos w=2u l=1u
M8415 n3910 n3838 VDD VDD pmos w=2u l=1u
M8416 n3910 n3838 VSS VSS nmos w=1u l=1u
M8417 n3832 n3913 VSS VSS nmos w=1u l=1u
M8418 n3832 n3912 VSS VSS nmos w=1u l=1u
M8419 n3832 n3913 net2537 VDD pmos w=2u l=1u
M8420 net2537 n3912 VDD VDD pmos w=2u l=1u
M8421 n3913 net2538 VSS VSS nmos w=1u l=1u
M8422 net2539 n3829 VSS VSS nmos w=1u l=1u
M8423 net2538 n3830 net2539 VSS nmos w=1u l=1u
M8424 net2538 n3829 VDD VDD pmos w=2u l=1u
M8425 net2538 n3830 VDD VDD pmos w=2u l=1u
M8426 n3913 net2538 VDD VDD pmos w=2u l=1u
M8427 n3912 n3828 VDD VDD pmos w=2u l=1u
M8428 n3912 n3828 VSS VSS nmos w=1u l=1u
M8429 n3822 n3915 VSS VSS nmos w=1u l=1u
M8430 n3822 n3914 VSS VSS nmos w=1u l=1u
M8431 n3822 n3915 net2540 VDD pmos w=2u l=1u
M8432 net2540 n3914 VDD VDD pmos w=2u l=1u
M8433 n3915 net2541 VSS VSS nmos w=1u l=1u
M8434 net2542 n3819 VSS VSS nmos w=1u l=1u
M8435 net2541 n3820 net2542 VSS nmos w=1u l=1u
M8436 net2541 n3819 VDD VDD pmos w=2u l=1u
M8437 net2541 n3820 VDD VDD pmos w=2u l=1u
M8438 n3915 net2541 VDD VDD pmos w=2u l=1u
M8439 n3914 n3818 VDD VDD pmos w=2u l=1u
M8440 n3914 n3818 VSS VSS nmos w=1u l=1u
M8441 n3812 n3917 VSS VSS nmos w=1u l=1u
M8442 n3812 n3916 VSS VSS nmos w=1u l=1u
M8443 n3812 n3917 net2543 VDD pmos w=2u l=1u
M8444 net2543 n3916 VDD VDD pmos w=2u l=1u
M8445 n3917 net2544 VSS VSS nmos w=1u l=1u
M8446 net2545 n3809 VSS VSS nmos w=1u l=1u
M8447 net2544 n3810 net2545 VSS nmos w=1u l=1u
M8448 net2544 n3809 VDD VDD pmos w=2u l=1u
M8449 net2544 n3810 VDD VDD pmos w=2u l=1u
M8450 n3917 net2544 VDD VDD pmos w=2u l=1u
M8451 n3916 n3808 VDD VDD pmos w=2u l=1u
M8452 n3916 n3808 VSS VSS nmos w=1u l=1u
M8453 n3802 n3919 VSS VSS nmos w=1u l=1u
M8454 n3802 n3918 VSS VSS nmos w=1u l=1u
M8455 n3802 n3919 net2546 VDD pmos w=2u l=1u
M8456 net2546 n3918 VDD VDD pmos w=2u l=1u
M8457 n3919 n3921 VSS VSS nmos w=1u l=1u
M8458 n3919 n3920 VSS VSS nmos w=1u l=1u
M8459 n3919 n3921 net2547 VDD pmos w=2u l=1u
M8460 net2547 n3920 VDD VDD pmos w=2u l=1u
M8461 n3920 n3800 VDD VDD pmos w=2u l=1u
M8462 n3920 n3800 VSS VSS nmos w=1u l=1u
M8463 n3918 n3798 VDD VDD pmos w=2u l=1u
M8464 n3918 n3798 VSS VSS nmos w=1u l=1u
M8465 n3791 n3923 VSS VSS nmos w=1u l=1u
M8466 n3791 n3922 VSS VSS nmos w=1u l=1u
M8467 n3791 n3923 net2548 VDD pmos w=2u l=1u
M8468 net2548 n3922 VDD VDD pmos w=2u l=1u
M8469 n3923 n3925 VSS VSS nmos w=1u l=1u
M8470 n3923 n3924 VSS VSS nmos w=1u l=1u
M8471 n3923 n3925 net2549 VDD pmos w=2u l=1u
M8472 net2549 n3924 VDD VDD pmos w=2u l=1u
M8473 n3924 n3790 VDD VDD pmos w=2u l=1u
M8474 n3924 n3790 VSS VSS nmos w=1u l=1u
M8475 n3922 n3788 VDD VDD pmos w=2u l=1u
M8476 n3922 n3788 VSS VSS nmos w=1u l=1u
M8477 n3781 n3927 VSS VSS nmos w=1u l=1u
M8478 n3781 n3926 VSS VSS nmos w=1u l=1u
M8479 n3781 n3927 net2550 VDD pmos w=2u l=1u
M8480 net2550 n3926 VDD VDD pmos w=2u l=1u
M8481 n3927 n3779 VSS VSS nmos w=1u l=1u
M8482 n3927 n3780 VSS VSS nmos w=1u l=1u
M8483 n3927 n3779 net2551 VDD pmos w=2u l=1u
M8484 net2551 n3780 VDD VDD pmos w=2u l=1u
M8485 n3926 n3778 VDD VDD pmos w=2u l=1u
M8486 n3926 n3778 VSS VSS nmos w=1u l=1u
M8487 net2552 n3780 VSS VSS nmos w=1u l=1u
M8488 net2553 n3928 VSS VSS nmos w=1u l=1u
M8489 N5672 net2554 VSS VSS nmos w=1u l=1u
M8490 net2554 n3780 net2555 VSS nmos w=1u l=1u
M8491 net2554 net2552 net2553 VSS nmos w=1u l=1u
M8492 net2555 net2553 VSS VSS nmos w=1u l=1u
M8493 net2554 net2552 net2556 VDD pmos w=2u l=1u
M8494 net2552 n3780 VDD VDD pmos w=2u l=1u
M8495 net2553 n3780 net2554 VDD pmos w=2u l=1u
M8496 net2553 n3928 VDD VDD pmos w=2u l=1u
M8497 N5672 net2554 VDD VDD pmos w=2u l=1u
M8498 net2556 net2553 VDD VDD pmos w=2u l=1u
M8499 n3780 n2271 VSS VSS nmos w=1u l=1u
M8500 n3780 n3929 VSS VSS nmos w=1u l=1u
M8501 n3780 n2271 net2557 VDD pmos w=2u l=1u
M8502 net2557 n3929 VDD VDD pmos w=2u l=1u
M8503 n2271 N494 VDD VDD pmos w=2u l=1u
M8504 n2271 N494 VSS VSS nmos w=1u l=1u
M8505 n3928 n3779 VDD VDD pmos w=2u l=1u
M8506 n3928 n3779 VSS VSS nmos w=1u l=1u
M8507 n3779 n3778 net2558 VSS nmos w=1u l=1u
M8508 net2558 n3930 VSS VSS nmos w=1u l=1u
M8509 n3779 n3778 VDD VDD pmos w=2u l=1u
M8510 n3779 n3930 VDD VDD pmos w=2u l=1u
M8511 n3778 n3932 net2559 VSS nmos w=1u l=1u
M8512 net2559 n3931 VSS VSS nmos w=1u l=1u
M8513 n3778 n3932 VDD VDD pmos w=2u l=1u
M8514 n3778 n3931 VDD VDD pmos w=2u l=1u
M8515 n3932 n3934 net2560 VSS nmos w=1u l=1u
M8516 net2560 n3933 VSS VSS nmos w=1u l=1u
M8517 n3932 n3934 VDD VDD pmos w=2u l=1u
M8518 n3932 n3933 VDD VDD pmos w=2u l=1u
M8519 n3933 net2561 VSS VSS nmos w=1u l=1u
M8520 net2561 n3935 VSS VSS nmos w=1u l=1u
M8521 net2561 n3936 VSS VSS nmos w=1u l=1u
M8522 net2561 n3936 net2562 VDD pmos w=2u l=1u
M8523 n3933 net2561 VDD VDD pmos w=2u l=1u
M8524 net2562 n3935 VDD VDD pmos w=2u l=1u
M8525 net2563 n3789 VSS VSS nmos w=1u l=1u
M8526 net2564 n3790 VSS VSS nmos w=1u l=1u
M8527 n3931 net2565 VSS VSS nmos w=1u l=1u
M8528 net2565 n3789 net2566 VSS nmos w=1u l=1u
M8529 net2565 net2563 net2564 VSS nmos w=1u l=1u
M8530 net2566 net2564 VSS VSS nmos w=1u l=1u
M8531 net2565 net2563 net2567 VDD pmos w=2u l=1u
M8532 net2563 n3789 VDD VDD pmos w=2u l=1u
M8533 net2564 n3789 net2565 VDD pmos w=2u l=1u
M8534 net2564 n3790 VDD VDD pmos w=2u l=1u
M8535 n3931 net2565 VDD VDD pmos w=2u l=1u
M8536 net2567 net2564 VDD VDD pmos w=2u l=1u
M8537 n3789 n3925 VDD VDD pmos w=2u l=1u
M8538 n3789 n3925 VSS VSS nmos w=1u l=1u
M8539 n3930 n3938 net2568 VSS nmos w=1u l=1u
M8540 net2568 n3937 VSS VSS nmos w=1u l=1u
M8541 n3930 n3938 VDD VDD pmos w=2u l=1u
M8542 n3930 n3937 VDD VDD pmos w=2u l=1u
M8543 net2569 n3790 VSS VSS nmos w=1u l=1u
M8544 net2570 n3925 VSS VSS nmos w=1u l=1u
M8545 n3938 net2571 VSS VSS nmos w=1u l=1u
M8546 net2571 n3790 net2572 VSS nmos w=1u l=1u
M8547 net2571 net2569 net2570 VSS nmos w=1u l=1u
M8548 net2572 net2570 VSS VSS nmos w=1u l=1u
M8549 net2571 net2569 net2573 VDD pmos w=2u l=1u
M8550 net2569 n3790 VDD VDD pmos w=2u l=1u
M8551 net2570 n3790 net2571 VDD pmos w=2u l=1u
M8552 net2570 n3925 VDD VDD pmos w=2u l=1u
M8553 n3938 net2571 VDD VDD pmos w=2u l=1u
M8554 net2573 net2570 VDD VDD pmos w=2u l=1u
M8555 n3790 N477 net2574 VSS nmos w=1u l=1u
M8556 net2574 N18 VSS VSS nmos w=1u l=1u
M8557 n3790 N477 VDD VDD pmos w=2u l=1u
M8558 n3790 N18 VDD VDD pmos w=2u l=1u
M8559 n3925 n3788 net2575 VSS nmos w=1u l=1u
M8560 net2575 n3939 VSS VSS nmos w=1u l=1u
M8561 n3925 n3788 VDD VDD pmos w=2u l=1u
M8562 n3925 n3939 VDD VDD pmos w=2u l=1u
M8563 n3788 n3941 net2576 VSS nmos w=1u l=1u
M8564 net2576 n3940 VSS VSS nmos w=1u l=1u
M8565 n3788 n3941 VDD VDD pmos w=2u l=1u
M8566 n3788 n3940 VDD VDD pmos w=2u l=1u
M8567 n3941 n3943 net2577 VSS nmos w=1u l=1u
M8568 net2577 n3942 VSS VSS nmos w=1u l=1u
M8569 n3941 n3943 VDD VDD pmos w=2u l=1u
M8570 n3941 n3942 VDD VDD pmos w=2u l=1u
M8571 n3942 n3945 net2578 VSS nmos w=1u l=1u
M8572 net2578 n3944 VSS VSS nmos w=1u l=1u
M8573 n3942 n3945 VDD VDD pmos w=2u l=1u
M8574 n3942 n3944 VDD VDD pmos w=2u l=1u
M8575 net2579 n3799 VSS VSS nmos w=1u l=1u
M8576 net2580 n3800 VSS VSS nmos w=1u l=1u
M8577 n3940 net2581 VSS VSS nmos w=1u l=1u
M8578 net2581 n3799 net2582 VSS nmos w=1u l=1u
M8579 net2581 net2579 net2580 VSS nmos w=1u l=1u
M8580 net2582 net2580 VSS VSS nmos w=1u l=1u
M8581 net2581 net2579 net2583 VDD pmos w=2u l=1u
M8582 net2579 n3799 VDD VDD pmos w=2u l=1u
M8583 net2580 n3799 net2581 VDD pmos w=2u l=1u
M8584 net2580 n3800 VDD VDD pmos w=2u l=1u
M8585 n3940 net2581 VDD VDD pmos w=2u l=1u
M8586 net2583 net2580 VDD VDD pmos w=2u l=1u
M8587 n3799 n3921 VDD VDD pmos w=2u l=1u
M8588 n3799 n3921 VSS VSS nmos w=1u l=1u
M8589 n3939 n3947 net2584 VSS nmos w=1u l=1u
M8590 net2584 n3946 VSS VSS nmos w=1u l=1u
M8591 n3939 n3947 VDD VDD pmos w=2u l=1u
M8592 n3939 n3946 VDD VDD pmos w=2u l=1u
M8593 net2585 n3800 VSS VSS nmos w=1u l=1u
M8594 net2586 n3921 VSS VSS nmos w=1u l=1u
M8595 n3947 net2587 VSS VSS nmos w=1u l=1u
M8596 net2587 n3800 net2588 VSS nmos w=1u l=1u
M8597 net2587 net2585 net2586 VSS nmos w=1u l=1u
M8598 net2588 net2586 VSS VSS nmos w=1u l=1u
M8599 net2587 net2585 net2589 VDD pmos w=2u l=1u
M8600 net2585 n3800 VDD VDD pmos w=2u l=1u
M8601 net2586 n3800 net2587 VDD pmos w=2u l=1u
M8602 net2586 n3921 VDD VDD pmos w=2u l=1u
M8603 n3947 net2587 VDD VDD pmos w=2u l=1u
M8604 net2589 net2586 VDD VDD pmos w=2u l=1u
M8605 n3800 N460 net2590 VSS nmos w=1u l=1u
M8606 net2590 N35 VSS VSS nmos w=1u l=1u
M8607 n3800 N460 VDD VDD pmos w=2u l=1u
M8608 n3800 N35 VDD VDD pmos w=2u l=1u
M8609 n3921 n3798 net2591 VSS nmos w=1u l=1u
M8610 net2591 n3948 VSS VSS nmos w=1u l=1u
M8611 n3921 n3798 VDD VDD pmos w=2u l=1u
M8612 n3921 n3948 VDD VDD pmos w=2u l=1u
M8613 n3798 n3950 net2592 VSS nmos w=1u l=1u
M8614 net2592 n3949 VSS VSS nmos w=1u l=1u
M8615 n3798 n3950 VDD VDD pmos w=2u l=1u
M8616 n3798 n3949 VDD VDD pmos w=2u l=1u
M8617 n3950 n3952 net2593 VSS nmos w=1u l=1u
M8618 net2593 n3951 VSS VSS nmos w=1u l=1u
M8619 n3950 n3952 VDD VDD pmos w=2u l=1u
M8620 n3950 n3951 VDD VDD pmos w=2u l=1u
M8621 n3951 n3954 net2594 VSS nmos w=1u l=1u
M8622 net2594 n3953 VSS VSS nmos w=1u l=1u
M8623 n3951 n3954 VDD VDD pmos w=2u l=1u
M8624 n3951 n3953 VDD VDD pmos w=2u l=1u
M8625 net2595 n3809 VSS VSS nmos w=1u l=1u
M8626 net2596 n3810 VSS VSS nmos w=1u l=1u
M8627 n3949 net2597 VSS VSS nmos w=1u l=1u
M8628 net2597 n3809 net2598 VSS nmos w=1u l=1u
M8629 net2597 net2595 net2596 VSS nmos w=1u l=1u
M8630 net2598 net2596 VSS VSS nmos w=1u l=1u
M8631 net2597 net2595 net2599 VDD pmos w=2u l=1u
M8632 net2595 n3809 VDD VDD pmos w=2u l=1u
M8633 net2596 n3809 net2597 VDD pmos w=2u l=1u
M8634 net2596 n3810 VDD VDD pmos w=2u l=1u
M8635 n3949 net2597 VDD VDD pmos w=2u l=1u
M8636 net2599 net2596 VDD VDD pmos w=2u l=1u
M8637 n3809 n3955 VDD VDD pmos w=2u l=1u
M8638 n3809 n3955 VSS VSS nmos w=1u l=1u
M8639 n3948 n3957 net2600 VSS nmos w=1u l=1u
M8640 net2600 n3956 VSS VSS nmos w=1u l=1u
M8641 n3948 n3957 VDD VDD pmos w=2u l=1u
M8642 n3948 n3956 VDD VDD pmos w=2u l=1u
M8643 net2601 n3810 VSS VSS nmos w=1u l=1u
M8644 net2602 n3955 VSS VSS nmos w=1u l=1u
M8645 n3957 net2603 VSS VSS nmos w=1u l=1u
M8646 net2603 n3810 net2604 VSS nmos w=1u l=1u
M8647 net2603 net2601 net2602 VSS nmos w=1u l=1u
M8648 net2604 net2602 VSS VSS nmos w=1u l=1u
M8649 net2603 net2601 net2605 VDD pmos w=2u l=1u
M8650 net2601 n3810 VDD VDD pmos w=2u l=1u
M8651 net2602 n3810 net2603 VDD pmos w=2u l=1u
M8652 net2602 n3955 VDD VDD pmos w=2u l=1u
M8653 n3957 net2603 VDD VDD pmos w=2u l=1u
M8654 net2605 net2602 VDD VDD pmos w=2u l=1u
M8655 n3810 N443 net2606 VSS nmos w=1u l=1u
M8656 net2606 N52 VSS VSS nmos w=1u l=1u
M8657 n3810 N443 VDD VDD pmos w=2u l=1u
M8658 n3810 N52 VDD VDD pmos w=2u l=1u
M8659 n3955 n3808 net2607 VSS nmos w=1u l=1u
M8660 net2607 n3958 VSS VSS nmos w=1u l=1u
M8661 n3955 n3808 VDD VDD pmos w=2u l=1u
M8662 n3955 n3958 VDD VDD pmos w=2u l=1u
M8663 n3808 n3960 net2608 VSS nmos w=1u l=1u
M8664 net2608 n3959 VSS VSS nmos w=1u l=1u
M8665 n3808 n3960 VDD VDD pmos w=2u l=1u
M8666 n3808 n3959 VDD VDD pmos w=2u l=1u
M8667 n3960 n3962 net2609 VSS nmos w=1u l=1u
M8668 net2609 n3961 VSS VSS nmos w=1u l=1u
M8669 n3960 n3962 VDD VDD pmos w=2u l=1u
M8670 n3960 n3961 VDD VDD pmos w=2u l=1u
M8671 n3961 n3964 net2610 VSS nmos w=1u l=1u
M8672 net2610 n3963 VSS VSS nmos w=1u l=1u
M8673 n3961 n3964 VDD VDD pmos w=2u l=1u
M8674 n3961 n3963 VDD VDD pmos w=2u l=1u
M8675 net2611 n3819 VSS VSS nmos w=1u l=1u
M8676 net2612 n3820 VSS VSS nmos w=1u l=1u
M8677 n3959 net2613 VSS VSS nmos w=1u l=1u
M8678 net2613 n3819 net2614 VSS nmos w=1u l=1u
M8679 net2613 net2611 net2612 VSS nmos w=1u l=1u
M8680 net2614 net2612 VSS VSS nmos w=1u l=1u
M8681 net2613 net2611 net2615 VDD pmos w=2u l=1u
M8682 net2611 n3819 VDD VDD pmos w=2u l=1u
M8683 net2612 n3819 net2613 VDD pmos w=2u l=1u
M8684 net2612 n3820 VDD VDD pmos w=2u l=1u
M8685 n3959 net2613 VDD VDD pmos w=2u l=1u
M8686 net2615 net2612 VDD VDD pmos w=2u l=1u
M8687 n3819 n3965 VDD VDD pmos w=2u l=1u
M8688 n3819 n3965 VSS VSS nmos w=1u l=1u
M8689 n3958 n3967 net2616 VSS nmos w=1u l=1u
M8690 net2616 n3966 VSS VSS nmos w=1u l=1u
M8691 n3958 n3967 VDD VDD pmos w=2u l=1u
M8692 n3958 n3966 VDD VDD pmos w=2u l=1u
M8693 net2617 n3820 VSS VSS nmos w=1u l=1u
M8694 net2618 n3965 VSS VSS nmos w=1u l=1u
M8695 n3967 net2619 VSS VSS nmos w=1u l=1u
M8696 net2619 n3820 net2620 VSS nmos w=1u l=1u
M8697 net2619 net2617 net2618 VSS nmos w=1u l=1u
M8698 net2620 net2618 VSS VSS nmos w=1u l=1u
M8699 net2619 net2617 net2621 VDD pmos w=2u l=1u
M8700 net2617 n3820 VDD VDD pmos w=2u l=1u
M8701 net2618 n3820 net2619 VDD pmos w=2u l=1u
M8702 net2618 n3965 VDD VDD pmos w=2u l=1u
M8703 n3967 net2619 VDD VDD pmos w=2u l=1u
M8704 net2621 net2618 VDD VDD pmos w=2u l=1u
M8705 n3820 N426 net2622 VSS nmos w=1u l=1u
M8706 net2622 N69 VSS VSS nmos w=1u l=1u
M8707 n3820 N426 VDD VDD pmos w=2u l=1u
M8708 n3820 N69 VDD VDD pmos w=2u l=1u
M8709 n3965 n3818 net2623 VSS nmos w=1u l=1u
M8710 net2623 n3968 VSS VSS nmos w=1u l=1u
M8711 n3965 n3818 VDD VDD pmos w=2u l=1u
M8712 n3965 n3968 VDD VDD pmos w=2u l=1u
M8713 n3818 n3970 net2624 VSS nmos w=1u l=1u
M8714 net2624 n3969 VSS VSS nmos w=1u l=1u
M8715 n3818 n3970 VDD VDD pmos w=2u l=1u
M8716 n3818 n3969 VDD VDD pmos w=2u l=1u
M8717 n3970 n3972 net2625 VSS nmos w=1u l=1u
M8718 net2625 n3971 VSS VSS nmos w=1u l=1u
M8719 n3970 n3972 VDD VDD pmos w=2u l=1u
M8720 n3970 n3971 VDD VDD pmos w=2u l=1u
M8721 n3971 n3974 net2626 VSS nmos w=1u l=1u
M8722 net2626 n3973 VSS VSS nmos w=1u l=1u
M8723 n3971 n3974 VDD VDD pmos w=2u l=1u
M8724 n3971 n3973 VDD VDD pmos w=2u l=1u
M8725 net2627 n3829 VSS VSS nmos w=1u l=1u
M8726 net2628 n3830 VSS VSS nmos w=1u l=1u
M8727 n3969 net2629 VSS VSS nmos w=1u l=1u
M8728 net2629 n3829 net2630 VSS nmos w=1u l=1u
M8729 net2629 net2627 net2628 VSS nmos w=1u l=1u
M8730 net2630 net2628 VSS VSS nmos w=1u l=1u
M8731 net2629 net2627 net2631 VDD pmos w=2u l=1u
M8732 net2627 n3829 VDD VDD pmos w=2u l=1u
M8733 net2628 n3829 net2629 VDD pmos w=2u l=1u
M8734 net2628 n3830 VDD VDD pmos w=2u l=1u
M8735 n3969 net2629 VDD VDD pmos w=2u l=1u
M8736 net2631 net2628 VDD VDD pmos w=2u l=1u
M8737 n3829 n3975 VDD VDD pmos w=2u l=1u
M8738 n3829 n3975 VSS VSS nmos w=1u l=1u
M8739 n3968 n3977 net2632 VSS nmos w=1u l=1u
M8740 net2632 n3976 VSS VSS nmos w=1u l=1u
M8741 n3968 n3977 VDD VDD pmos w=2u l=1u
M8742 n3968 n3976 VDD VDD pmos w=2u l=1u
M8743 net2633 n3830 VSS VSS nmos w=1u l=1u
M8744 net2634 n3975 VSS VSS nmos w=1u l=1u
M8745 n3977 net2635 VSS VSS nmos w=1u l=1u
M8746 net2635 n3830 net2636 VSS nmos w=1u l=1u
M8747 net2635 net2633 net2634 VSS nmos w=1u l=1u
M8748 net2636 net2634 VSS VSS nmos w=1u l=1u
M8749 net2635 net2633 net2637 VDD pmos w=2u l=1u
M8750 net2633 n3830 VDD VDD pmos w=2u l=1u
M8751 net2634 n3830 net2635 VDD pmos w=2u l=1u
M8752 net2634 n3975 VDD VDD pmos w=2u l=1u
M8753 n3977 net2635 VDD VDD pmos w=2u l=1u
M8754 net2637 net2634 VDD VDD pmos w=2u l=1u
M8755 n3830 N409 net2638 VSS nmos w=1u l=1u
M8756 net2638 N86 VSS VSS nmos w=1u l=1u
M8757 n3830 N409 VDD VDD pmos w=2u l=1u
M8758 n3830 N86 VDD VDD pmos w=2u l=1u
M8759 n3975 n3828 net2639 VSS nmos w=1u l=1u
M8760 net2639 n3978 VSS VSS nmos w=1u l=1u
M8761 n3975 n3828 VDD VDD pmos w=2u l=1u
M8762 n3975 n3978 VDD VDD pmos w=2u l=1u
M8763 n3828 n3980 net2640 VSS nmos w=1u l=1u
M8764 net2640 n3979 VSS VSS nmos w=1u l=1u
M8765 n3828 n3980 VDD VDD pmos w=2u l=1u
M8766 n3828 n3979 VDD VDD pmos w=2u l=1u
M8767 n3980 n3982 net2641 VSS nmos w=1u l=1u
M8768 net2641 n3981 VSS VSS nmos w=1u l=1u
M8769 n3980 n3982 VDD VDD pmos w=2u l=1u
M8770 n3980 n3981 VDD VDD pmos w=2u l=1u
M8771 n3981 n3984 net2642 VSS nmos w=1u l=1u
M8772 net2642 n3983 VSS VSS nmos w=1u l=1u
M8773 n3981 n3984 VDD VDD pmos w=2u l=1u
M8774 n3981 n3983 VDD VDD pmos w=2u l=1u
M8775 net2643 n3839 VSS VSS nmos w=1u l=1u
M8776 net2644 n3840 VSS VSS nmos w=1u l=1u
M8777 n3979 net2645 VSS VSS nmos w=1u l=1u
M8778 net2645 n3839 net2646 VSS nmos w=1u l=1u
M8779 net2645 net2643 net2644 VSS nmos w=1u l=1u
M8780 net2646 net2644 VSS VSS nmos w=1u l=1u
M8781 net2645 net2643 net2647 VDD pmos w=2u l=1u
M8782 net2643 n3839 VDD VDD pmos w=2u l=1u
M8783 net2644 n3839 net2645 VDD pmos w=2u l=1u
M8784 net2644 n3840 VDD VDD pmos w=2u l=1u
M8785 n3979 net2645 VDD VDD pmos w=2u l=1u
M8786 net2647 net2644 VDD VDD pmos w=2u l=1u
M8787 n3839 n3985 VDD VDD pmos w=2u l=1u
M8788 n3839 n3985 VSS VSS nmos w=1u l=1u
M8789 n3978 n3987 net2648 VSS nmos w=1u l=1u
M8790 net2648 n3986 VSS VSS nmos w=1u l=1u
M8791 n3978 n3987 VDD VDD pmos w=2u l=1u
M8792 n3978 n3986 VDD VDD pmos w=2u l=1u
M8793 net2649 n3840 VSS VSS nmos w=1u l=1u
M8794 net2650 n3985 VSS VSS nmos w=1u l=1u
M8795 n3987 net2651 VSS VSS nmos w=1u l=1u
M8796 net2651 n3840 net2652 VSS nmos w=1u l=1u
M8797 net2651 net2649 net2650 VSS nmos w=1u l=1u
M8798 net2652 net2650 VSS VSS nmos w=1u l=1u
M8799 net2651 net2649 net2653 VDD pmos w=2u l=1u
M8800 net2649 n3840 VDD VDD pmos w=2u l=1u
M8801 net2650 n3840 net2651 VDD pmos w=2u l=1u
M8802 net2650 n3985 VDD VDD pmos w=2u l=1u
M8803 n3987 net2651 VDD VDD pmos w=2u l=1u
M8804 net2653 net2650 VDD VDD pmos w=2u l=1u
M8805 n3840 N392 net2654 VSS nmos w=1u l=1u
M8806 net2654 N103 VSS VSS nmos w=1u l=1u
M8807 n3840 N392 VDD VDD pmos w=2u l=1u
M8808 n3840 N103 VDD VDD pmos w=2u l=1u
M8809 n3985 n3838 net2655 VSS nmos w=1u l=1u
M8810 net2655 n3988 VSS VSS nmos w=1u l=1u
M8811 n3985 n3838 VDD VDD pmos w=2u l=1u
M8812 n3985 n3988 VDD VDD pmos w=2u l=1u
M8813 n3838 n3990 net2656 VSS nmos w=1u l=1u
M8814 net2656 n3989 VSS VSS nmos w=1u l=1u
M8815 n3838 n3990 VDD VDD pmos w=2u l=1u
M8816 n3838 n3989 VDD VDD pmos w=2u l=1u
M8817 n3990 n3992 net2657 VSS nmos w=1u l=1u
M8818 net2657 n3991 VSS VSS nmos w=1u l=1u
M8819 n3990 n3992 VDD VDD pmos w=2u l=1u
M8820 n3990 n3991 VDD VDD pmos w=2u l=1u
M8821 n3991 n3994 net2658 VSS nmos w=1u l=1u
M8822 net2658 n3993 VSS VSS nmos w=1u l=1u
M8823 n3991 n3994 VDD VDD pmos w=2u l=1u
M8824 n3991 n3993 VDD VDD pmos w=2u l=1u
M8825 net2659 n3849 VSS VSS nmos w=1u l=1u
M8826 net2660 n3850 VSS VSS nmos w=1u l=1u
M8827 n3989 net2661 VSS VSS nmos w=1u l=1u
M8828 net2661 n3849 net2662 VSS nmos w=1u l=1u
M8829 net2661 net2659 net2660 VSS nmos w=1u l=1u
M8830 net2662 net2660 VSS VSS nmos w=1u l=1u
M8831 net2661 net2659 net2663 VDD pmos w=2u l=1u
M8832 net2659 n3849 VDD VDD pmos w=2u l=1u
M8833 net2660 n3849 net2661 VDD pmos w=2u l=1u
M8834 net2660 n3850 VDD VDD pmos w=2u l=1u
M8835 n3989 net2661 VDD VDD pmos w=2u l=1u
M8836 net2663 net2660 VDD VDD pmos w=2u l=1u
M8837 n3849 n3995 VDD VDD pmos w=2u l=1u
M8838 n3849 n3995 VSS VSS nmos w=1u l=1u
M8839 n3988 n3997 net2664 VSS nmos w=1u l=1u
M8840 net2664 n3996 VSS VSS nmos w=1u l=1u
M8841 n3988 n3997 VDD VDD pmos w=2u l=1u
M8842 n3988 n3996 VDD VDD pmos w=2u l=1u
M8843 net2665 n3850 VSS VSS nmos w=1u l=1u
M8844 net2666 n3995 VSS VSS nmos w=1u l=1u
M8845 n3997 net2667 VSS VSS nmos w=1u l=1u
M8846 net2667 n3850 net2668 VSS nmos w=1u l=1u
M8847 net2667 net2665 net2666 VSS nmos w=1u l=1u
M8848 net2668 net2666 VSS VSS nmos w=1u l=1u
M8849 net2667 net2665 net2669 VDD pmos w=2u l=1u
M8850 net2665 n3850 VDD VDD pmos w=2u l=1u
M8851 net2666 n3850 net2667 VDD pmos w=2u l=1u
M8852 net2666 n3995 VDD VDD pmos w=2u l=1u
M8853 n3997 net2667 VDD VDD pmos w=2u l=1u
M8854 net2669 net2666 VDD VDD pmos w=2u l=1u
M8855 n3850 N375 net2670 VSS nmos w=1u l=1u
M8856 net2670 N120 VSS VSS nmos w=1u l=1u
M8857 n3850 N375 VDD VDD pmos w=2u l=1u
M8858 n3850 N120 VDD VDD pmos w=2u l=1u
M8859 n3995 n3848 net2671 VSS nmos w=1u l=1u
M8860 net2671 n3998 VSS VSS nmos w=1u l=1u
M8861 n3995 n3848 VDD VDD pmos w=2u l=1u
M8862 n3995 n3998 VDD VDD pmos w=2u l=1u
M8863 n3848 n4000 net2672 VSS nmos w=1u l=1u
M8864 net2672 n3999 VSS VSS nmos w=1u l=1u
M8865 n3848 n4000 VDD VDD pmos w=2u l=1u
M8866 n3848 n3999 VDD VDD pmos w=2u l=1u
M8867 n4000 n4002 net2673 VSS nmos w=1u l=1u
M8868 net2673 n4001 VSS VSS nmos w=1u l=1u
M8869 n4000 n4002 VDD VDD pmos w=2u l=1u
M8870 n4000 n4001 VDD VDD pmos w=2u l=1u
M8871 n4001 net2674 VSS VSS nmos w=1u l=1u
M8872 net2674 n4003 VSS VSS nmos w=1u l=1u
M8873 net2674 n4004 VSS VSS nmos w=1u l=1u
M8874 net2674 n4004 net2675 VDD pmos w=2u l=1u
M8875 n4001 net2674 VDD VDD pmos w=2u l=1u
M8876 net2675 n4003 VDD VDD pmos w=2u l=1u
M8877 net2676 n3859 VSS VSS nmos w=1u l=1u
M8878 net2677 n3860 VSS VSS nmos w=1u l=1u
M8879 n3999 net2678 VSS VSS nmos w=1u l=1u
M8880 net2678 n3859 net2679 VSS nmos w=1u l=1u
M8881 net2678 net2676 net2677 VSS nmos w=1u l=1u
M8882 net2679 net2677 VSS VSS nmos w=1u l=1u
M8883 net2678 net2676 net2680 VDD pmos w=2u l=1u
M8884 net2676 n3859 VDD VDD pmos w=2u l=1u
M8885 net2677 n3859 net2678 VDD pmos w=2u l=1u
M8886 net2677 n3860 VDD VDD pmos w=2u l=1u
M8887 n3999 net2678 VDD VDD pmos w=2u l=1u
M8888 net2680 net2677 VDD VDD pmos w=2u l=1u
M8889 n3860 n4005 VDD VDD pmos w=2u l=1u
M8890 n3860 n4005 VSS VSS nmos w=1u l=1u
M8891 n3998 n4007 net2681 VSS nmos w=1u l=1u
M8892 net2681 n4006 VSS VSS nmos w=1u l=1u
M8893 n3998 n4007 VDD VDD pmos w=2u l=1u
M8894 n3998 n4006 VDD VDD pmos w=2u l=1u
M8895 net2682 n4005 VSS VSS nmos w=1u l=1u
M8896 net2683 n3859 VSS VSS nmos w=1u l=1u
M8897 n4007 net2684 VSS VSS nmos w=1u l=1u
M8898 net2684 n4005 net2685 VSS nmos w=1u l=1u
M8899 net2684 net2682 net2683 VSS nmos w=1u l=1u
M8900 net2685 net2683 VSS VSS nmos w=1u l=1u
M8901 net2684 net2682 net2686 VDD pmos w=2u l=1u
M8902 net2682 n4005 VDD VDD pmos w=2u l=1u
M8903 net2683 n4005 net2684 VDD pmos w=2u l=1u
M8904 net2683 n3859 VDD VDD pmos w=2u l=1u
M8905 n4007 net2684 VDD VDD pmos w=2u l=1u
M8906 net2686 net2683 VDD VDD pmos w=2u l=1u
M8907 n4005 N358 net2687 VSS nmos w=1u l=1u
M8908 net2687 N137 VSS VSS nmos w=1u l=1u
M8909 n4005 N358 VDD VDD pmos w=2u l=1u
M8910 n4005 N137 VDD VDD pmos w=2u l=1u
M8911 n3859 n3858 net2688 VSS nmos w=1u l=1u
M8912 net2688 n4008 VSS VSS nmos w=1u l=1u
M8913 n3859 n3858 VDD VDD pmos w=2u l=1u
M8914 n3859 n4008 VDD VDD pmos w=2u l=1u
M8915 n3858 n4010 net2689 VSS nmos w=1u l=1u
M8916 net2689 n4009 VSS VSS nmos w=1u l=1u
M8917 n3858 n4010 VDD VDD pmos w=2u l=1u
M8918 n3858 n4009 VDD VDD pmos w=2u l=1u
M8919 n4010 n4012 net2690 VSS nmos w=1u l=1u
M8920 net2690 n4011 VSS VSS nmos w=1u l=1u
M8921 n4010 n4012 VDD VDD pmos w=2u l=1u
M8922 n4010 n4011 VDD VDD pmos w=2u l=1u
M8923 n4011 n4014 net2691 VSS nmos w=1u l=1u
M8924 net2691 n4013 VSS VSS nmos w=1u l=1u
M8925 n4011 n4014 VDD VDD pmos w=2u l=1u
M8926 n4011 n4013 VDD VDD pmos w=2u l=1u
M8927 net2692 n3869 VSS VSS nmos w=1u l=1u
M8928 net2693 n3870 VSS VSS nmos w=1u l=1u
M8929 n4009 net2694 VSS VSS nmos w=1u l=1u
M8930 net2694 n3869 net2695 VSS nmos w=1u l=1u
M8931 net2694 net2692 net2693 VSS nmos w=1u l=1u
M8932 net2695 net2693 VSS VSS nmos w=1u l=1u
M8933 net2694 net2692 net2696 VDD pmos w=2u l=1u
M8934 net2692 n3869 VDD VDD pmos w=2u l=1u
M8935 net2693 n3869 net2694 VDD pmos w=2u l=1u
M8936 net2693 n3870 VDD VDD pmos w=2u l=1u
M8937 n4009 net2694 VDD VDD pmos w=2u l=1u
M8938 net2696 net2693 VDD VDD pmos w=2u l=1u
M8939 n3869 n4015 VDD VDD pmos w=2u l=1u
M8940 n3869 n4015 VSS VSS nmos w=1u l=1u
M8941 n4008 n4017 net2697 VSS nmos w=1u l=1u
M8942 net2697 n4016 VSS VSS nmos w=1u l=1u
M8943 n4008 n4017 VDD VDD pmos w=2u l=1u
M8944 n4008 n4016 VDD VDD pmos w=2u l=1u
M8945 net2698 n3870 VSS VSS nmos w=1u l=1u
M8946 net2699 n4015 VSS VSS nmos w=1u l=1u
M8947 n4017 net2700 VSS VSS nmos w=1u l=1u
M8948 net2700 n3870 net2701 VSS nmos w=1u l=1u
M8949 net2700 net2698 net2699 VSS nmos w=1u l=1u
M8950 net2701 net2699 VSS VSS nmos w=1u l=1u
M8951 net2700 net2698 net2702 VDD pmos w=2u l=1u
M8952 net2698 n3870 VDD VDD pmos w=2u l=1u
M8953 net2699 n3870 net2700 VDD pmos w=2u l=1u
M8954 net2699 n4015 VDD VDD pmos w=2u l=1u
M8955 n4017 net2700 VDD VDD pmos w=2u l=1u
M8956 net2702 net2699 VDD VDD pmos w=2u l=1u
M8957 n3870 N341 net2703 VSS nmos w=1u l=1u
M8958 net2703 N154 VSS VSS nmos w=1u l=1u
M8959 n3870 N341 VDD VDD pmos w=2u l=1u
M8960 n3870 N154 VDD VDD pmos w=2u l=1u
M8961 n4015 n3868 net2704 VSS nmos w=1u l=1u
M8962 net2704 n4018 VSS VSS nmos w=1u l=1u
M8963 n4015 n3868 VDD VDD pmos w=2u l=1u
M8964 n4015 n4018 VDD VDD pmos w=2u l=1u
M8965 n3868 n4020 net2705 VSS nmos w=1u l=1u
M8966 net2705 n4019 VSS VSS nmos w=1u l=1u
M8967 n3868 n4020 VDD VDD pmos w=2u l=1u
M8968 n3868 n4019 VDD VDD pmos w=2u l=1u
M8969 n4020 net2706 VSS VSS nmos w=1u l=1u
M8970 net2706 n4021 VSS VSS nmos w=1u l=1u
M8971 net2706 n4022 VSS VSS nmos w=1u l=1u
M8972 net2706 n4022 net2707 VDD pmos w=2u l=1u
M8973 n4020 net2706 VDD VDD pmos w=2u l=1u
M8974 net2707 n4021 VDD VDD pmos w=2u l=1u
M8975 n4019 net2708 VSS VSS nmos w=1u l=1u
M8976 net2709 n4023 VSS VSS nmos w=1u l=1u
M8977 net2708 n3903 net2709 VSS nmos w=1u l=1u
M8978 net2708 n4023 VDD VDD pmos w=2u l=1u
M8979 net2708 n3903 VDD VDD pmos w=2u l=1u
M8980 n4019 net2708 VDD VDD pmos w=2u l=1u
M8981 n4018 n4025 net2710 VSS nmos w=1u l=1u
M8982 net2710 n4024 VSS VSS nmos w=1u l=1u
M8983 n4018 n4025 VDD VDD pmos w=2u l=1u
M8984 n4018 n4024 VDD VDD pmos w=2u l=1u
M8985 n4025 n3903 net2711 VSS nmos w=1u l=1u
M8986 net2711 n4023 VSS VSS nmos w=1u l=1u
M8987 n4025 n3903 VDD VDD pmos w=2u l=1u
M8988 n4025 n4023 VDD VDD pmos w=2u l=1u
M8989 n3903 n4027 net2712 VSS nmos w=1u l=1u
M8990 net2712 n4026 VSS VSS nmos w=1u l=1u
M8991 n3903 n4027 VDD VDD pmos w=2u l=1u
M8992 n3903 n4026 VDD VDD pmos w=2u l=1u
M8993 n4027 N324 net2713 VSS nmos w=1u l=1u
M8994 net2713 N171 VSS VSS nmos w=1u l=1u
M8995 n4027 N324 VDD VDD pmos w=2u l=1u
M8996 n4027 N171 VDD VDD pmos w=2u l=1u
M8997 n4023 N171 net2714 VSS nmos w=1u l=1u
M8998 net2714 n4028 VSS VSS nmos w=1u l=1u
M8999 n4023 N171 VDD VDD pmos w=2u l=1u
M9000 n4023 n4028 VDD VDD pmos w=2u l=1u
M9001 n4028 n3257 VSS VSS nmos w=1u l=1u
M9002 n4028 n4026 VSS VSS nmos w=1u l=1u
M9003 n4028 n3257 net2715 VDD pmos w=2u l=1u
M9004 net2715 n4026 VDD VDD pmos w=2u l=1u
M9005 n4026 n3878 VSS VSS nmos w=1u l=1u
M9006 n4026 n4029 VSS VSS nmos w=1u l=1u
M9007 n4026 n3878 net2716 VDD pmos w=2u l=1u
M9008 net2716 n4029 VDD VDD pmos w=2u l=1u
M9009 n3878 n4031 VSS VSS nmos w=1u l=1u
M9010 n3878 n4030 VSS VSS nmos w=1u l=1u
M9011 n3878 n4031 net2717 VDD pmos w=2u l=1u
M9012 net2717 n4030 VDD VDD pmos w=2u l=1u
M9013 n4029 net2718 VSS VSS nmos w=1u l=1u
M9014 net2719 n4030 VSS VSS nmos w=1u l=1u
M9015 net2718 n4031 net2719 VSS nmos w=1u l=1u
M9016 net2718 n4030 VDD VDD pmos w=2u l=1u
M9017 net2718 n4031 VDD VDD pmos w=2u l=1u
M9018 n4029 net2718 VDD VDD pmos w=2u l=1u
M9019 n4030 n4032 net2720 VSS nmos w=1u l=1u
M9020 net2720 n3901 VSS VSS nmos w=1u l=1u
M9021 n4030 n4032 VDD VDD pmos w=2u l=1u
M9022 n4030 n3901 VDD VDD pmos w=2u l=1u
M9023 n4032 N188 net2721 VSS nmos w=1u l=1u
M9024 net2721 n4033 VSS VSS nmos w=1u l=1u
M9025 n4032 N188 VDD VDD pmos w=2u l=1u
M9026 n4032 n4033 VDD VDD pmos w=2u l=1u
M9027 n4033 n3411 VSS VSS nmos w=1u l=1u
M9028 n4033 n4034 VSS VSS nmos w=1u l=1u
M9029 n4033 n3411 net2722 VDD pmos w=2u l=1u
M9030 net2722 n4034 VDD VDD pmos w=2u l=1u
M9031 n3901 n4035 net2723 VSS nmos w=1u l=1u
M9032 net2723 n4034 VSS VSS nmos w=1u l=1u
M9033 n3901 n4035 VDD VDD pmos w=2u l=1u
M9034 n3901 n4034 VDD VDD pmos w=2u l=1u
M9035 n4035 N307 net2724 VSS nmos w=1u l=1u
M9036 net2724 N188 VSS VSS nmos w=1u l=1u
M9037 n4035 N307 VDD VDD pmos w=2u l=1u
M9038 n4035 N188 VDD VDD pmos w=2u l=1u
M9039 n4034 net2725 VSS VSS nmos w=1u l=1u
M9040 net2726 n4036 VSS VSS nmos w=1u l=1u
M9041 net2725 n3902 net2726 VSS nmos w=1u l=1u
M9042 net2725 n4036 VDD VDD pmos w=2u l=1u
M9043 net2725 n3902 VDD VDD pmos w=2u l=1u
M9044 n4034 net2725 VDD VDD pmos w=2u l=1u
M9045 n4036 n3893 net2727 VSS nmos w=1u l=1u
M9046 net2727 n4037 VSS VSS nmos w=1u l=1u
M9047 n4036 n3893 VDD VDD pmos w=2u l=1u
M9048 n4036 n4037 VDD VDD pmos w=2u l=1u
M9049 n3902 n4039 net2728 VSS nmos w=1u l=1u
M9050 net2728 n4038 VSS VSS nmos w=1u l=1u
M9051 n3902 n4039 VDD VDD pmos w=2u l=1u
M9052 n3902 n4038 VDD VDD pmos w=2u l=1u
M9053 n4039 n3893 net2729 VSS nmos w=1u l=1u
M9054 net2729 n4040 VSS VSS nmos w=1u l=1u
M9055 n4039 n3893 VDD VDD pmos w=2u l=1u
M9056 n4039 n4040 VDD VDD pmos w=2u l=1u
M9057 n3893 N205 net2730 VSS nmos w=1u l=1u
M9058 net2730 n4041 VSS VSS nmos w=1u l=1u
M9059 n3893 N205 VDD VDD pmos w=2u l=1u
M9060 n3893 n4041 VDD VDD pmos w=2u l=1u
M9061 n4041 net2731 VSS VSS nmos w=1u l=1u
M9062 net2732 N222 VSS VSS nmos w=1u l=1u
M9063 net2731 n3741 net2732 VSS nmos w=1u l=1u
M9064 net2731 N222 VDD VDD pmos w=2u l=1u
M9065 net2731 n3741 VDD VDD pmos w=2u l=1u
M9066 n4041 net2731 VDD VDD pmos w=2u l=1u
M9067 n4040 n4043 net2733 VSS nmos w=1u l=1u
M9068 net2733 n4042 VSS VSS nmos w=1u l=1u
M9069 n4040 n4043 VDD VDD pmos w=2u l=1u
M9070 n4040 n4042 VDD VDD pmos w=2u l=1u
M9071 n4043 N273 net2734 VSS nmos w=1u l=1u
M9072 net2734 N222 VSS VSS nmos w=1u l=1u
M9073 n4043 N273 VDD VDD pmos w=2u l=1u
M9074 n4043 N222 VDD VDD pmos w=2u l=1u
M9075 n4042 N290 net2735 VSS nmos w=1u l=1u
M9076 net2735 N205 VSS VSS nmos w=1u l=1u
M9077 n4042 N290 VDD VDD pmos w=2u l=1u
M9078 n4042 N205 VDD VDD pmos w=2u l=1u
M9079 n4031 net2736 VSS VSS nmos w=1u l=1u
M9080 net2737 n4045 VSS VSS nmos w=1u l=1u
M9081 net2736 n4044 net2737 VSS nmos w=1u l=1u
M9082 net2736 n4045 VDD VDD pmos w=2u l=1u
M9083 net2736 n4044 VDD VDD pmos w=2u l=1u
M9084 n4031 net2736 VDD VDD pmos w=2u l=1u
M9085 n4024 n4021 VSS VSS nmos w=1u l=1u
M9086 n4024 n4022 VSS VSS nmos w=1u l=1u
M9087 n4024 n4021 net2738 VDD pmos w=2u l=1u
M9088 net2738 n4022 VDD VDD pmos w=2u l=1u
M9089 n4021 n4046 VDD VDD pmos w=2u l=1u
M9090 n4021 n4046 VSS VSS nmos w=1u l=1u
M9091 n4016 n4048 VSS VSS nmos w=1u l=1u
M9092 n4016 n4047 VSS VSS nmos w=1u l=1u
M9093 n4016 n4048 net2739 VDD pmos w=2u l=1u
M9094 net2739 n4047 VDD VDD pmos w=2u l=1u
M9095 n4048 net2740 VSS VSS nmos w=1u l=1u
M9096 net2741 n4013 VSS VSS nmos w=1u l=1u
M9097 net2740 n4014 net2741 VSS nmos w=1u l=1u
M9098 net2740 n4013 VDD VDD pmos w=2u l=1u
M9099 net2740 n4014 VDD VDD pmos w=2u l=1u
M9100 n4048 net2740 VDD VDD pmos w=2u l=1u
M9101 n4047 n4012 VDD VDD pmos w=2u l=1u
M9102 n4047 n4012 VSS VSS nmos w=1u l=1u
M9103 n4006 n4050 VSS VSS nmos w=1u l=1u
M9104 n4006 n4049 VSS VSS nmos w=1u l=1u
M9105 n4006 n4050 net2742 VDD pmos w=2u l=1u
M9106 net2742 n4049 VDD VDD pmos w=2u l=1u
M9107 n4050 n4003 VSS VSS nmos w=1u l=1u
M9108 n4050 n4004 VSS VSS nmos w=1u l=1u
M9109 n4050 n4003 net2743 VDD pmos w=2u l=1u
M9110 net2743 n4004 VDD VDD pmos w=2u l=1u
M9111 n4049 n4002 VDD VDD pmos w=2u l=1u
M9112 n4049 n4002 VSS VSS nmos w=1u l=1u
M9113 n3996 n4052 VSS VSS nmos w=1u l=1u
M9114 n3996 n4051 VSS VSS nmos w=1u l=1u
M9115 n3996 n4052 net2744 VDD pmos w=2u l=1u
M9116 net2744 n4051 VDD VDD pmos w=2u l=1u
M9117 n4052 net2745 VSS VSS nmos w=1u l=1u
M9118 net2746 n3993 VSS VSS nmos w=1u l=1u
M9119 net2745 n3994 net2746 VSS nmos w=1u l=1u
M9120 net2745 n3993 VDD VDD pmos w=2u l=1u
M9121 net2745 n3994 VDD VDD pmos w=2u l=1u
M9122 n4052 net2745 VDD VDD pmos w=2u l=1u
M9123 n4051 n3992 VDD VDD pmos w=2u l=1u
M9124 n4051 n3992 VSS VSS nmos w=1u l=1u
M9125 n3986 n4054 VSS VSS nmos w=1u l=1u
M9126 n3986 n4053 VSS VSS nmos w=1u l=1u
M9127 n3986 n4054 net2747 VDD pmos w=2u l=1u
M9128 net2747 n4053 VDD VDD pmos w=2u l=1u
M9129 n4054 net2748 VSS VSS nmos w=1u l=1u
M9130 net2749 n3983 VSS VSS nmos w=1u l=1u
M9131 net2748 n3984 net2749 VSS nmos w=1u l=1u
M9132 net2748 n3983 VDD VDD pmos w=2u l=1u
M9133 net2748 n3984 VDD VDD pmos w=2u l=1u
M9134 n4054 net2748 VDD VDD pmos w=2u l=1u
M9135 n4053 n3982 VDD VDD pmos w=2u l=1u
M9136 n4053 n3982 VSS VSS nmos w=1u l=1u
M9137 n3976 n4056 VSS VSS nmos w=1u l=1u
M9138 n3976 n4055 VSS VSS nmos w=1u l=1u
M9139 n3976 n4056 net2750 VDD pmos w=2u l=1u
M9140 net2750 n4055 VDD VDD pmos w=2u l=1u
M9141 n4056 net2751 VSS VSS nmos w=1u l=1u
M9142 net2752 n3973 VSS VSS nmos w=1u l=1u
M9143 net2751 n3974 net2752 VSS nmos w=1u l=1u
M9144 net2751 n3973 VDD VDD pmos w=2u l=1u
M9145 net2751 n3974 VDD VDD pmos w=2u l=1u
M9146 n4056 net2751 VDD VDD pmos w=2u l=1u
M9147 n4055 n3972 VDD VDD pmos w=2u l=1u
M9148 n4055 n3972 VSS VSS nmos w=1u l=1u
M9149 n3966 n4058 VSS VSS nmos w=1u l=1u
M9150 n3966 n4057 VSS VSS nmos w=1u l=1u
M9151 n3966 n4058 net2753 VDD pmos w=2u l=1u
M9152 net2753 n4057 VDD VDD pmos w=2u l=1u
M9153 n4058 net2754 VSS VSS nmos w=1u l=1u
M9154 net2755 n3963 VSS VSS nmos w=1u l=1u
M9155 net2754 n3964 net2755 VSS nmos w=1u l=1u
M9156 net2754 n3963 VDD VDD pmos w=2u l=1u
M9157 net2754 n3964 VDD VDD pmos w=2u l=1u
M9158 n4058 net2754 VDD VDD pmos w=2u l=1u
M9159 n4057 n3962 VDD VDD pmos w=2u l=1u
M9160 n4057 n3962 VSS VSS nmos w=1u l=1u
M9161 n3956 n4060 VSS VSS nmos w=1u l=1u
M9162 n3956 n4059 VSS VSS nmos w=1u l=1u
M9163 n3956 n4060 net2756 VDD pmos w=2u l=1u
M9164 net2756 n4059 VDD VDD pmos w=2u l=1u
M9165 n4060 n4062 VSS VSS nmos w=1u l=1u
M9166 n4060 n4061 VSS VSS nmos w=1u l=1u
M9167 n4060 n4062 net2757 VDD pmos w=2u l=1u
M9168 net2757 n4061 VDD VDD pmos w=2u l=1u
M9169 n4061 n3954 VDD VDD pmos w=2u l=1u
M9170 n4061 n3954 VSS VSS nmos w=1u l=1u
M9171 n4059 n3952 VDD VDD pmos w=2u l=1u
M9172 n4059 n3952 VSS VSS nmos w=1u l=1u
M9173 n3946 n4064 VSS VSS nmos w=1u l=1u
M9174 n3946 n4063 VSS VSS nmos w=1u l=1u
M9175 n3946 n4064 net2758 VDD pmos w=2u l=1u
M9176 net2758 n4063 VDD VDD pmos w=2u l=1u
M9177 n4064 n4066 VSS VSS nmos w=1u l=1u
M9178 n4064 n4065 VSS VSS nmos w=1u l=1u
M9179 n4064 n4066 net2759 VDD pmos w=2u l=1u
M9180 net2759 n4065 VDD VDD pmos w=2u l=1u
M9181 n4065 n3945 VDD VDD pmos w=2u l=1u
M9182 n4065 n3945 VSS VSS nmos w=1u l=1u
M9183 n4063 n3943 VDD VDD pmos w=2u l=1u
M9184 n4063 n3943 VSS VSS nmos w=1u l=1u
M9185 n3937 n4068 VSS VSS nmos w=1u l=1u
M9186 n3937 n4067 VSS VSS nmos w=1u l=1u
M9187 n3937 n4068 net2760 VDD pmos w=2u l=1u
M9188 net2760 n4067 VDD VDD pmos w=2u l=1u
M9189 n4068 n3935 VSS VSS nmos w=1u l=1u
M9190 n4068 n3936 VSS VSS nmos w=1u l=1u
M9191 n4068 n3935 net2761 VDD pmos w=2u l=1u
M9192 net2761 n3936 VDD VDD pmos w=2u l=1u
M9193 n4067 n3934 VDD VDD pmos w=2u l=1u
M9194 n4067 n3934 VSS VSS nmos w=1u l=1u
M9195 net2762 n3936 VSS VSS nmos w=1u l=1u
M9196 net2763 n4069 VSS VSS nmos w=1u l=1u
M9197 N5308 net2764 VSS VSS nmos w=1u l=1u
M9198 net2764 n3936 net2765 VSS nmos w=1u l=1u
M9199 net2764 net2762 net2763 VSS nmos w=1u l=1u
M9200 net2765 net2763 VSS VSS nmos w=1u l=1u
M9201 net2764 net2762 net2766 VDD pmos w=2u l=1u
M9202 net2762 n3936 VDD VDD pmos w=2u l=1u
M9203 net2763 n3936 net2764 VDD pmos w=2u l=1u
M9204 net2763 n4069 VDD VDD pmos w=2u l=1u
M9205 N5308 net2764 VDD VDD pmos w=2u l=1u
M9206 net2766 net2763 VDD VDD pmos w=2u l=1u
M9207 n3936 n2321 VSS VSS nmos w=1u l=1u
M9208 n3936 n3929 VSS VSS nmos w=1u l=1u
M9209 n3936 n2321 net2767 VDD pmos w=2u l=1u
M9210 net2767 n3929 VDD VDD pmos w=2u l=1u
M9211 n2321 N477 VDD VDD pmos w=2u l=1u
M9212 n2321 N477 VSS VSS nmos w=1u l=1u
M9213 n4069 n3935 VDD VDD pmos w=2u l=1u
M9214 n4069 n3935 VSS VSS nmos w=1u l=1u
M9215 n3935 n3934 net2768 VSS nmos w=1u l=1u
M9216 net2768 n4070 VSS VSS nmos w=1u l=1u
M9217 n3935 n3934 VDD VDD pmos w=2u l=1u
M9218 n3935 n4070 VDD VDD pmos w=2u l=1u
M9219 n3934 n4072 net2769 VSS nmos w=1u l=1u
M9220 net2769 n4071 VSS VSS nmos w=1u l=1u
M9221 n3934 n4072 VDD VDD pmos w=2u l=1u
M9222 n3934 n4071 VDD VDD pmos w=2u l=1u
M9223 n4072 n4074 net2770 VSS nmos w=1u l=1u
M9224 net2770 n4073 VSS VSS nmos w=1u l=1u
M9225 n4072 n4074 VDD VDD pmos w=2u l=1u
M9226 n4072 n4073 VDD VDD pmos w=2u l=1u
M9227 n4073 net2771 VSS VSS nmos w=1u l=1u
M9228 net2771 n4075 VSS VSS nmos w=1u l=1u
M9229 net2771 n4076 VSS VSS nmos w=1u l=1u
M9230 net2771 n4076 net2772 VDD pmos w=2u l=1u
M9231 n4073 net2771 VDD VDD pmos w=2u l=1u
M9232 net2772 n4075 VDD VDD pmos w=2u l=1u
M9233 net2773 n3944 VSS VSS nmos w=1u l=1u
M9234 net2774 n3945 VSS VSS nmos w=1u l=1u
M9235 n4071 net2775 VSS VSS nmos w=1u l=1u
M9236 net2775 n3944 net2776 VSS nmos w=1u l=1u
M9237 net2775 net2773 net2774 VSS nmos w=1u l=1u
M9238 net2776 net2774 VSS VSS nmos w=1u l=1u
M9239 net2775 net2773 net2777 VDD pmos w=2u l=1u
M9240 net2773 n3944 VDD VDD pmos w=2u l=1u
M9241 net2774 n3944 net2775 VDD pmos w=2u l=1u
M9242 net2774 n3945 VDD VDD pmos w=2u l=1u
M9243 n4071 net2775 VDD VDD pmos w=2u l=1u
M9244 net2777 net2774 VDD VDD pmos w=2u l=1u
M9245 n3944 n4066 VDD VDD pmos w=2u l=1u
M9246 n3944 n4066 VSS VSS nmos w=1u l=1u
M9247 n4070 n4078 net2778 VSS nmos w=1u l=1u
M9248 net2778 n4077 VSS VSS nmos w=1u l=1u
M9249 n4070 n4078 VDD VDD pmos w=2u l=1u
M9250 n4070 n4077 VDD VDD pmos w=2u l=1u
M9251 net2779 n3945 VSS VSS nmos w=1u l=1u
M9252 net2780 n4066 VSS VSS nmos w=1u l=1u
M9253 n4078 net2781 VSS VSS nmos w=1u l=1u
M9254 net2781 n3945 net2782 VSS nmos w=1u l=1u
M9255 net2781 net2779 net2780 VSS nmos w=1u l=1u
M9256 net2782 net2780 VSS VSS nmos w=1u l=1u
M9257 net2781 net2779 net2783 VDD pmos w=2u l=1u
M9258 net2779 n3945 VDD VDD pmos w=2u l=1u
M9259 net2780 n3945 net2781 VDD pmos w=2u l=1u
M9260 net2780 n4066 VDD VDD pmos w=2u l=1u
M9261 n4078 net2781 VDD VDD pmos w=2u l=1u
M9262 net2783 net2780 VDD VDD pmos w=2u l=1u
M9263 n3945 N460 net2784 VSS nmos w=1u l=1u
M9264 net2784 N18 VSS VSS nmos w=1u l=1u
M9265 n3945 N460 VDD VDD pmos w=2u l=1u
M9266 n3945 N18 VDD VDD pmos w=2u l=1u
M9267 n4066 n3943 net2785 VSS nmos w=1u l=1u
M9268 net2785 n4079 VSS VSS nmos w=1u l=1u
M9269 n4066 n3943 VDD VDD pmos w=2u l=1u
M9270 n4066 n4079 VDD VDD pmos w=2u l=1u
M9271 n3943 n4081 net2786 VSS nmos w=1u l=1u
M9272 net2786 n4080 VSS VSS nmos w=1u l=1u
M9273 n3943 n4081 VDD VDD pmos w=2u l=1u
M9274 n3943 n4080 VDD VDD pmos w=2u l=1u
M9275 n4081 n4083 net2787 VSS nmos w=1u l=1u
M9276 net2787 n4082 VSS VSS nmos w=1u l=1u
M9277 n4081 n4083 VDD VDD pmos w=2u l=1u
M9278 n4081 n4082 VDD VDD pmos w=2u l=1u
M9279 n4082 n4085 net2788 VSS nmos w=1u l=1u
M9280 net2788 n4084 VSS VSS nmos w=1u l=1u
M9281 n4082 n4085 VDD VDD pmos w=2u l=1u
M9282 n4082 n4084 VDD VDD pmos w=2u l=1u
M9283 net2789 n3953 VSS VSS nmos w=1u l=1u
M9284 net2790 n3954 VSS VSS nmos w=1u l=1u
M9285 n4080 net2791 VSS VSS nmos w=1u l=1u
M9286 net2791 n3953 net2792 VSS nmos w=1u l=1u
M9287 net2791 net2789 net2790 VSS nmos w=1u l=1u
M9288 net2792 net2790 VSS VSS nmos w=1u l=1u
M9289 net2791 net2789 net2793 VDD pmos w=2u l=1u
M9290 net2789 n3953 VDD VDD pmos w=2u l=1u
M9291 net2790 n3953 net2791 VDD pmos w=2u l=1u
M9292 net2790 n3954 VDD VDD pmos w=2u l=1u
M9293 n4080 net2791 VDD VDD pmos w=2u l=1u
M9294 net2793 net2790 VDD VDD pmos w=2u l=1u
M9295 n3953 n4062 VDD VDD pmos w=2u l=1u
M9296 n3953 n4062 VSS VSS nmos w=1u l=1u
M9297 n4079 n4087 net2794 VSS nmos w=1u l=1u
M9298 net2794 n4086 VSS VSS nmos w=1u l=1u
M9299 n4079 n4087 VDD VDD pmos w=2u l=1u
M9300 n4079 n4086 VDD VDD pmos w=2u l=1u
M9301 net2795 n3954 VSS VSS nmos w=1u l=1u
M9302 net2796 n4062 VSS VSS nmos w=1u l=1u
M9303 n4087 net2797 VSS VSS nmos w=1u l=1u
M9304 net2797 n3954 net2798 VSS nmos w=1u l=1u
M9305 net2797 net2795 net2796 VSS nmos w=1u l=1u
M9306 net2798 net2796 VSS VSS nmos w=1u l=1u
M9307 net2797 net2795 net2799 VDD pmos w=2u l=1u
M9308 net2795 n3954 VDD VDD pmos w=2u l=1u
M9309 net2796 n3954 net2797 VDD pmos w=2u l=1u
M9310 net2796 n4062 VDD VDD pmos w=2u l=1u
M9311 n4087 net2797 VDD VDD pmos w=2u l=1u
M9312 net2799 net2796 VDD VDD pmos w=2u l=1u
M9313 n3954 N443 net2800 VSS nmos w=1u l=1u
M9314 net2800 N35 VSS VSS nmos w=1u l=1u
M9315 n3954 N443 VDD VDD pmos w=2u l=1u
M9316 n3954 N35 VDD VDD pmos w=2u l=1u
M9317 n4062 n3952 net2801 VSS nmos w=1u l=1u
M9318 net2801 n4088 VSS VSS nmos w=1u l=1u
M9319 n4062 n3952 VDD VDD pmos w=2u l=1u
M9320 n4062 n4088 VDD VDD pmos w=2u l=1u
M9321 n3952 n4090 net2802 VSS nmos w=1u l=1u
M9322 net2802 n4089 VSS VSS nmos w=1u l=1u
M9323 n3952 n4090 VDD VDD pmos w=2u l=1u
M9324 n3952 n4089 VDD VDD pmos w=2u l=1u
M9325 n4090 n4092 net2803 VSS nmos w=1u l=1u
M9326 net2803 n4091 VSS VSS nmos w=1u l=1u
M9327 n4090 n4092 VDD VDD pmos w=2u l=1u
M9328 n4090 n4091 VDD VDD pmos w=2u l=1u
M9329 n4091 n4094 net2804 VSS nmos w=1u l=1u
M9330 net2804 n4093 VSS VSS nmos w=1u l=1u
M9331 n4091 n4094 VDD VDD pmos w=2u l=1u
M9332 n4091 n4093 VDD VDD pmos w=2u l=1u
M9333 net2805 n3963 VSS VSS nmos w=1u l=1u
M9334 net2806 n3964 VSS VSS nmos w=1u l=1u
M9335 n4089 net2807 VSS VSS nmos w=1u l=1u
M9336 net2807 n3963 net2808 VSS nmos w=1u l=1u
M9337 net2807 net2805 net2806 VSS nmos w=1u l=1u
M9338 net2808 net2806 VSS VSS nmos w=1u l=1u
M9339 net2807 net2805 net2809 VDD pmos w=2u l=1u
M9340 net2805 n3963 VDD VDD pmos w=2u l=1u
M9341 net2806 n3963 net2807 VDD pmos w=2u l=1u
M9342 net2806 n3964 VDD VDD pmos w=2u l=1u
M9343 n4089 net2807 VDD VDD pmos w=2u l=1u
M9344 net2809 net2806 VDD VDD pmos w=2u l=1u
M9345 n3963 n4095 VDD VDD pmos w=2u l=1u
M9346 n3963 n4095 VSS VSS nmos w=1u l=1u
M9347 n4088 n4097 net2810 VSS nmos w=1u l=1u
M9348 net2810 n4096 VSS VSS nmos w=1u l=1u
M9349 n4088 n4097 VDD VDD pmos w=2u l=1u
M9350 n4088 n4096 VDD VDD pmos w=2u l=1u
M9351 net2811 n3964 VSS VSS nmos w=1u l=1u
M9352 net2812 n4095 VSS VSS nmos w=1u l=1u
M9353 n4097 net2813 VSS VSS nmos w=1u l=1u
M9354 net2813 n3964 net2814 VSS nmos w=1u l=1u
M9355 net2813 net2811 net2812 VSS nmos w=1u l=1u
M9356 net2814 net2812 VSS VSS nmos w=1u l=1u
M9357 net2813 net2811 net2815 VDD pmos w=2u l=1u
M9358 net2811 n3964 VDD VDD pmos w=2u l=1u
M9359 net2812 n3964 net2813 VDD pmos w=2u l=1u
M9360 net2812 n4095 VDD VDD pmos w=2u l=1u
M9361 n4097 net2813 VDD VDD pmos w=2u l=1u
M9362 net2815 net2812 VDD VDD pmos w=2u l=1u
M9363 n3964 N426 net2816 VSS nmos w=1u l=1u
M9364 net2816 N52 VSS VSS nmos w=1u l=1u
M9365 n3964 N426 VDD VDD pmos w=2u l=1u
M9366 n3964 N52 VDD VDD pmos w=2u l=1u
M9367 n4095 n3962 net2817 VSS nmos w=1u l=1u
M9368 net2817 n4098 VSS VSS nmos w=1u l=1u
M9369 n4095 n3962 VDD VDD pmos w=2u l=1u
M9370 n4095 n4098 VDD VDD pmos w=2u l=1u
M9371 n3962 n4100 net2818 VSS nmos w=1u l=1u
M9372 net2818 n4099 VSS VSS nmos w=1u l=1u
M9373 n3962 n4100 VDD VDD pmos w=2u l=1u
M9374 n3962 n4099 VDD VDD pmos w=2u l=1u
M9375 n4100 n4102 net2819 VSS nmos w=1u l=1u
M9376 net2819 n4101 VSS VSS nmos w=1u l=1u
M9377 n4100 n4102 VDD VDD pmos w=2u l=1u
M9378 n4100 n4101 VDD VDD pmos w=2u l=1u
M9379 n4101 n4104 net2820 VSS nmos w=1u l=1u
M9380 net2820 n4103 VSS VSS nmos w=1u l=1u
M9381 n4101 n4104 VDD VDD pmos w=2u l=1u
M9382 n4101 n4103 VDD VDD pmos w=2u l=1u
M9383 net2821 n3973 VSS VSS nmos w=1u l=1u
M9384 net2822 n3974 VSS VSS nmos w=1u l=1u
M9385 n4099 net2823 VSS VSS nmos w=1u l=1u
M9386 net2823 n3973 net2824 VSS nmos w=1u l=1u
M9387 net2823 net2821 net2822 VSS nmos w=1u l=1u
M9388 net2824 net2822 VSS VSS nmos w=1u l=1u
M9389 net2823 net2821 net2825 VDD pmos w=2u l=1u
M9390 net2821 n3973 VDD VDD pmos w=2u l=1u
M9391 net2822 n3973 net2823 VDD pmos w=2u l=1u
M9392 net2822 n3974 VDD VDD pmos w=2u l=1u
M9393 n4099 net2823 VDD VDD pmos w=2u l=1u
M9394 net2825 net2822 VDD VDD pmos w=2u l=1u
M9395 n3973 n4105 VDD VDD pmos w=2u l=1u
M9396 n3973 n4105 VSS VSS nmos w=1u l=1u
M9397 n4098 n4107 net2826 VSS nmos w=1u l=1u
M9398 net2826 n4106 VSS VSS nmos w=1u l=1u
M9399 n4098 n4107 VDD VDD pmos w=2u l=1u
M9400 n4098 n4106 VDD VDD pmos w=2u l=1u
M9401 net2827 n3974 VSS VSS nmos w=1u l=1u
M9402 net2828 n4105 VSS VSS nmos w=1u l=1u
M9403 n4107 net2829 VSS VSS nmos w=1u l=1u
M9404 net2829 n3974 net2830 VSS nmos w=1u l=1u
M9405 net2829 net2827 net2828 VSS nmos w=1u l=1u
M9406 net2830 net2828 VSS VSS nmos w=1u l=1u
M9407 net2829 net2827 net2831 VDD pmos w=2u l=1u
M9408 net2827 n3974 VDD VDD pmos w=2u l=1u
M9409 net2828 n3974 net2829 VDD pmos w=2u l=1u
M9410 net2828 n4105 VDD VDD pmos w=2u l=1u
M9411 n4107 net2829 VDD VDD pmos w=2u l=1u
M9412 net2831 net2828 VDD VDD pmos w=2u l=1u
M9413 n3974 N409 net2832 VSS nmos w=1u l=1u
M9414 net2832 N69 VSS VSS nmos w=1u l=1u
M9415 n3974 N409 VDD VDD pmos w=2u l=1u
M9416 n3974 N69 VDD VDD pmos w=2u l=1u
M9417 n4105 n3972 net2833 VSS nmos w=1u l=1u
M9418 net2833 n4108 VSS VSS nmos w=1u l=1u
M9419 n4105 n3972 VDD VDD pmos w=2u l=1u
M9420 n4105 n4108 VDD VDD pmos w=2u l=1u
M9421 n3972 n4110 net2834 VSS nmos w=1u l=1u
M9422 net2834 n4109 VSS VSS nmos w=1u l=1u
M9423 n3972 n4110 VDD VDD pmos w=2u l=1u
M9424 n3972 n4109 VDD VDD pmos w=2u l=1u
M9425 n4110 n4112 net2835 VSS nmos w=1u l=1u
M9426 net2835 n4111 VSS VSS nmos w=1u l=1u
M9427 n4110 n4112 VDD VDD pmos w=2u l=1u
M9428 n4110 n4111 VDD VDD pmos w=2u l=1u
M9429 n4111 n4114 net2836 VSS nmos w=1u l=1u
M9430 net2836 n4113 VSS VSS nmos w=1u l=1u
M9431 n4111 n4114 VDD VDD pmos w=2u l=1u
M9432 n4111 n4113 VDD VDD pmos w=2u l=1u
M9433 net2837 n3983 VSS VSS nmos w=1u l=1u
M9434 net2838 n3984 VSS VSS nmos w=1u l=1u
M9435 n4109 net2839 VSS VSS nmos w=1u l=1u
M9436 net2839 n3983 net2840 VSS nmos w=1u l=1u
M9437 net2839 net2837 net2838 VSS nmos w=1u l=1u
M9438 net2840 net2838 VSS VSS nmos w=1u l=1u
M9439 net2839 net2837 net2841 VDD pmos w=2u l=1u
M9440 net2837 n3983 VDD VDD pmos w=2u l=1u
M9441 net2838 n3983 net2839 VDD pmos w=2u l=1u
M9442 net2838 n3984 VDD VDD pmos w=2u l=1u
M9443 n4109 net2839 VDD VDD pmos w=2u l=1u
M9444 net2841 net2838 VDD VDD pmos w=2u l=1u
M9445 n3983 n4115 VDD VDD pmos w=2u l=1u
M9446 n3983 n4115 VSS VSS nmos w=1u l=1u
M9447 n4108 n4117 net2842 VSS nmos w=1u l=1u
M9448 net2842 n4116 VSS VSS nmos w=1u l=1u
M9449 n4108 n4117 VDD VDD pmos w=2u l=1u
M9450 n4108 n4116 VDD VDD pmos w=2u l=1u
M9451 net2843 n3984 VSS VSS nmos w=1u l=1u
M9452 net2844 n4115 VSS VSS nmos w=1u l=1u
M9453 n4117 net2845 VSS VSS nmos w=1u l=1u
M9454 net2845 n3984 net2846 VSS nmos w=1u l=1u
M9455 net2845 net2843 net2844 VSS nmos w=1u l=1u
M9456 net2846 net2844 VSS VSS nmos w=1u l=1u
M9457 net2845 net2843 net2847 VDD pmos w=2u l=1u
M9458 net2843 n3984 VDD VDD pmos w=2u l=1u
M9459 net2844 n3984 net2845 VDD pmos w=2u l=1u
M9460 net2844 n4115 VDD VDD pmos w=2u l=1u
M9461 n4117 net2845 VDD VDD pmos w=2u l=1u
M9462 net2847 net2844 VDD VDD pmos w=2u l=1u
M9463 n3984 N392 net2848 VSS nmos w=1u l=1u
M9464 net2848 N86 VSS VSS nmos w=1u l=1u
M9465 n3984 N392 VDD VDD pmos w=2u l=1u
M9466 n3984 N86 VDD VDD pmos w=2u l=1u
M9467 n4115 n3982 net2849 VSS nmos w=1u l=1u
M9468 net2849 n4118 VSS VSS nmos w=1u l=1u
M9469 n4115 n3982 VDD VDD pmos w=2u l=1u
M9470 n4115 n4118 VDD VDD pmos w=2u l=1u
M9471 n3982 n4120 net2850 VSS nmos w=1u l=1u
M9472 net2850 n4119 VSS VSS nmos w=1u l=1u
M9473 n3982 n4120 VDD VDD pmos w=2u l=1u
M9474 n3982 n4119 VDD VDD pmos w=2u l=1u
M9475 n4120 n4122 net2851 VSS nmos w=1u l=1u
M9476 net2851 n4121 VSS VSS nmos w=1u l=1u
M9477 n4120 n4122 VDD VDD pmos w=2u l=1u
M9478 n4120 n4121 VDD VDD pmos w=2u l=1u
M9479 n4121 n4124 net2852 VSS nmos w=1u l=1u
M9480 net2852 n4123 VSS VSS nmos w=1u l=1u
M9481 n4121 n4124 VDD VDD pmos w=2u l=1u
M9482 n4121 n4123 VDD VDD pmos w=2u l=1u
M9483 net2853 n3993 VSS VSS nmos w=1u l=1u
M9484 net2854 n3994 VSS VSS nmos w=1u l=1u
M9485 n4119 net2855 VSS VSS nmos w=1u l=1u
M9486 net2855 n3993 net2856 VSS nmos w=1u l=1u
M9487 net2855 net2853 net2854 VSS nmos w=1u l=1u
M9488 net2856 net2854 VSS VSS nmos w=1u l=1u
M9489 net2855 net2853 net2857 VDD pmos w=2u l=1u
M9490 net2853 n3993 VDD VDD pmos w=2u l=1u
M9491 net2854 n3993 net2855 VDD pmos w=2u l=1u
M9492 net2854 n3994 VDD VDD pmos w=2u l=1u
M9493 n4119 net2855 VDD VDD pmos w=2u l=1u
M9494 net2857 net2854 VDD VDD pmos w=2u l=1u
M9495 n3993 n4125 VDD VDD pmos w=2u l=1u
M9496 n3993 n4125 VSS VSS nmos w=1u l=1u
M9497 n4118 n4127 net2858 VSS nmos w=1u l=1u
M9498 net2858 n4126 VSS VSS nmos w=1u l=1u
M9499 n4118 n4127 VDD VDD pmos w=2u l=1u
M9500 n4118 n4126 VDD VDD pmos w=2u l=1u
M9501 net2859 n3994 VSS VSS nmos w=1u l=1u
M9502 net2860 n4125 VSS VSS nmos w=1u l=1u
M9503 n4127 net2861 VSS VSS nmos w=1u l=1u
M9504 net2861 n3994 net2862 VSS nmos w=1u l=1u
M9505 net2861 net2859 net2860 VSS nmos w=1u l=1u
M9506 net2862 net2860 VSS VSS nmos w=1u l=1u
M9507 net2861 net2859 net2863 VDD pmos w=2u l=1u
M9508 net2859 n3994 VDD VDD pmos w=2u l=1u
M9509 net2860 n3994 net2861 VDD pmos w=2u l=1u
M9510 net2860 n4125 VDD VDD pmos w=2u l=1u
M9511 n4127 net2861 VDD VDD pmos w=2u l=1u
M9512 net2863 net2860 VDD VDD pmos w=2u l=1u
M9513 n3994 N375 net2864 VSS nmos w=1u l=1u
M9514 net2864 N103 VSS VSS nmos w=1u l=1u
M9515 n3994 N375 VDD VDD pmos w=2u l=1u
M9516 n3994 N103 VDD VDD pmos w=2u l=1u
M9517 n4125 n3992 net2865 VSS nmos w=1u l=1u
M9518 net2865 n4128 VSS VSS nmos w=1u l=1u
M9519 n4125 n3992 VDD VDD pmos w=2u l=1u
M9520 n4125 n4128 VDD VDD pmos w=2u l=1u
M9521 n3992 n4130 net2866 VSS nmos w=1u l=1u
M9522 net2866 n4129 VSS VSS nmos w=1u l=1u
M9523 n3992 n4130 VDD VDD pmos w=2u l=1u
M9524 n3992 n4129 VDD VDD pmos w=2u l=1u
M9525 n4130 n4132 net2867 VSS nmos w=1u l=1u
M9526 net2867 n4131 VSS VSS nmos w=1u l=1u
M9527 n4130 n4132 VDD VDD pmos w=2u l=1u
M9528 n4130 n4131 VDD VDD pmos w=2u l=1u
M9529 n4131 net2868 VSS VSS nmos w=1u l=1u
M9530 net2868 n4133 VSS VSS nmos w=1u l=1u
M9531 net2868 n4134 VSS VSS nmos w=1u l=1u
M9532 net2868 n4134 net2869 VDD pmos w=2u l=1u
M9533 n4131 net2868 VDD VDD pmos w=2u l=1u
M9534 net2869 n4133 VDD VDD pmos w=2u l=1u
M9535 net2870 n4003 VSS VSS nmos w=1u l=1u
M9536 net2871 n4004 VSS VSS nmos w=1u l=1u
M9537 n4129 net2872 VSS VSS nmos w=1u l=1u
M9538 net2872 n4003 net2873 VSS nmos w=1u l=1u
M9539 net2872 net2870 net2871 VSS nmos w=1u l=1u
M9540 net2873 net2871 VSS VSS nmos w=1u l=1u
M9541 net2872 net2870 net2874 VDD pmos w=2u l=1u
M9542 net2870 n4003 VDD VDD pmos w=2u l=1u
M9543 net2871 n4003 net2872 VDD pmos w=2u l=1u
M9544 net2871 n4004 VDD VDD pmos w=2u l=1u
M9545 n4129 net2872 VDD VDD pmos w=2u l=1u
M9546 net2874 net2871 VDD VDD pmos w=2u l=1u
M9547 n4004 n4135 VDD VDD pmos w=2u l=1u
M9548 n4004 n4135 VSS VSS nmos w=1u l=1u
M9549 n4128 n4137 net2875 VSS nmos w=1u l=1u
M9550 net2875 n4136 VSS VSS nmos w=1u l=1u
M9551 n4128 n4137 VDD VDD pmos w=2u l=1u
M9552 n4128 n4136 VDD VDD pmos w=2u l=1u
M9553 net2876 n4135 VSS VSS nmos w=1u l=1u
M9554 net2877 n4003 VSS VSS nmos w=1u l=1u
M9555 n4137 net2878 VSS VSS nmos w=1u l=1u
M9556 net2878 n4135 net2879 VSS nmos w=1u l=1u
M9557 net2878 net2876 net2877 VSS nmos w=1u l=1u
M9558 net2879 net2877 VSS VSS nmos w=1u l=1u
M9559 net2878 net2876 net2880 VDD pmos w=2u l=1u
M9560 net2876 n4135 VDD VDD pmos w=2u l=1u
M9561 net2877 n4135 net2878 VDD pmos w=2u l=1u
M9562 net2877 n4003 VDD VDD pmos w=2u l=1u
M9563 n4137 net2878 VDD VDD pmos w=2u l=1u
M9564 net2880 net2877 VDD VDD pmos w=2u l=1u
M9565 n4135 N358 net2881 VSS nmos w=1u l=1u
M9566 net2881 N120 VSS VSS nmos w=1u l=1u
M9567 n4135 N358 VDD VDD pmos w=2u l=1u
M9568 n4135 N120 VDD VDD pmos w=2u l=1u
M9569 n4003 n4002 net2882 VSS nmos w=1u l=1u
M9570 net2882 n4138 VSS VSS nmos w=1u l=1u
M9571 n4003 n4002 VDD VDD pmos w=2u l=1u
M9572 n4003 n4138 VDD VDD pmos w=2u l=1u
M9573 n4002 n4140 net2883 VSS nmos w=1u l=1u
M9574 net2883 n4139 VSS VSS nmos w=1u l=1u
M9575 n4002 n4140 VDD VDD pmos w=2u l=1u
M9576 n4002 n4139 VDD VDD pmos w=2u l=1u
M9577 n4140 n4142 net2884 VSS nmos w=1u l=1u
M9578 net2884 n4141 VSS VSS nmos w=1u l=1u
M9579 n4140 n4142 VDD VDD pmos w=2u l=1u
M9580 n4140 n4141 VDD VDD pmos w=2u l=1u
M9581 n4141 n4144 net2885 VSS nmos w=1u l=1u
M9582 net2885 n4143 VSS VSS nmos w=1u l=1u
M9583 n4141 n4144 VDD VDD pmos w=2u l=1u
M9584 n4141 n4143 VDD VDD pmos w=2u l=1u
M9585 net2886 n4013 VSS VSS nmos w=1u l=1u
M9586 net2887 n4014 VSS VSS nmos w=1u l=1u
M9587 n4139 net2888 VSS VSS nmos w=1u l=1u
M9588 net2888 n4013 net2889 VSS nmos w=1u l=1u
M9589 net2888 net2886 net2887 VSS nmos w=1u l=1u
M9590 net2889 net2887 VSS VSS nmos w=1u l=1u
M9591 net2888 net2886 net2890 VDD pmos w=2u l=1u
M9592 net2886 n4013 VDD VDD pmos w=2u l=1u
M9593 net2887 n4013 net2888 VDD pmos w=2u l=1u
M9594 net2887 n4014 VDD VDD pmos w=2u l=1u
M9595 n4139 net2888 VDD VDD pmos w=2u l=1u
M9596 net2890 net2887 VDD VDD pmos w=2u l=1u
M9597 n4013 n4145 VDD VDD pmos w=2u l=1u
M9598 n4013 n4145 VSS VSS nmos w=1u l=1u
M9599 n4138 n4147 net2891 VSS nmos w=1u l=1u
M9600 net2891 n4146 VSS VSS nmos w=1u l=1u
M9601 n4138 n4147 VDD VDD pmos w=2u l=1u
M9602 n4138 n4146 VDD VDD pmos w=2u l=1u
M9603 net2892 n4014 VSS VSS nmos w=1u l=1u
M9604 net2893 n4145 VSS VSS nmos w=1u l=1u
M9605 n4147 net2894 VSS VSS nmos w=1u l=1u
M9606 net2894 n4014 net2895 VSS nmos w=1u l=1u
M9607 net2894 net2892 net2893 VSS nmos w=1u l=1u
M9608 net2895 net2893 VSS VSS nmos w=1u l=1u
M9609 net2894 net2892 net2896 VDD pmos w=2u l=1u
M9610 net2892 n4014 VDD VDD pmos w=2u l=1u
M9611 net2893 n4014 net2894 VDD pmos w=2u l=1u
M9612 net2893 n4145 VDD VDD pmos w=2u l=1u
M9613 n4147 net2894 VDD VDD pmos w=2u l=1u
M9614 net2896 net2893 VDD VDD pmos w=2u l=1u
M9615 n4014 N341 net2897 VSS nmos w=1u l=1u
M9616 net2897 N137 VSS VSS nmos w=1u l=1u
M9617 n4014 N341 VDD VDD pmos w=2u l=1u
M9618 n4014 N137 VDD VDD pmos w=2u l=1u
M9619 n4145 n4012 net2898 VSS nmos w=1u l=1u
M9620 net2898 n4148 VSS VSS nmos w=1u l=1u
M9621 n4145 n4012 VDD VDD pmos w=2u l=1u
M9622 n4145 n4148 VDD VDD pmos w=2u l=1u
M9623 n4012 n4150 net2899 VSS nmos w=1u l=1u
M9624 net2899 n4149 VSS VSS nmos w=1u l=1u
M9625 n4012 n4150 VDD VDD pmos w=2u l=1u
M9626 n4012 n4149 VDD VDD pmos w=2u l=1u
M9627 n4150 net2900 VSS VSS nmos w=1u l=1u
M9628 net2900 n4151 VSS VSS nmos w=1u l=1u
M9629 net2900 n4152 VSS VSS nmos w=1u l=1u
M9630 net2900 n4152 net2901 VDD pmos w=2u l=1u
M9631 n4150 net2900 VDD VDD pmos w=2u l=1u
M9632 net2901 n4151 VDD VDD pmos w=2u l=1u
M9633 n4149 net2902 VSS VSS nmos w=1u l=1u
M9634 net2903 n4153 VSS VSS nmos w=1u l=1u
M9635 net2902 n4046 net2903 VSS nmos w=1u l=1u
M9636 net2902 n4153 VDD VDD pmos w=2u l=1u
M9637 net2902 n4046 VDD VDD pmos w=2u l=1u
M9638 n4149 net2902 VDD VDD pmos w=2u l=1u
M9639 n4148 n4155 net2904 VSS nmos w=1u l=1u
M9640 net2904 n4154 VSS VSS nmos w=1u l=1u
M9641 n4148 n4155 VDD VDD pmos w=2u l=1u
M9642 n4148 n4154 VDD VDD pmos w=2u l=1u
M9643 n4155 n4046 net2905 VSS nmos w=1u l=1u
M9644 net2905 n4153 VSS VSS nmos w=1u l=1u
M9645 n4155 n4046 VDD VDD pmos w=2u l=1u
M9646 n4155 n4153 VDD VDD pmos w=2u l=1u
M9647 n4046 n4157 net2906 VSS nmos w=1u l=1u
M9648 net2906 n4156 VSS VSS nmos w=1u l=1u
M9649 n4046 n4157 VDD VDD pmos w=2u l=1u
M9650 n4046 n4156 VDD VDD pmos w=2u l=1u
M9651 n4157 N324 net2907 VSS nmos w=1u l=1u
M9652 net2907 N154 VSS VSS nmos w=1u l=1u
M9653 n4157 N324 VDD VDD pmos w=2u l=1u
M9654 n4157 N154 VDD VDD pmos w=2u l=1u
M9655 n4153 N154 net2908 VSS nmos w=1u l=1u
M9656 net2908 n4158 VSS VSS nmos w=1u l=1u
M9657 n4153 N154 VDD VDD pmos w=2u l=1u
M9658 n4153 n4158 VDD VDD pmos w=2u l=1u
M9659 n4158 n3257 VSS VSS nmos w=1u l=1u
M9660 n4158 n4156 VSS VSS nmos w=1u l=1u
M9661 n4158 n3257 net2909 VDD pmos w=2u l=1u
M9662 net2909 n4156 VDD VDD pmos w=2u l=1u
M9663 n4156 n4022 VSS VSS nmos w=1u l=1u
M9664 n4156 n4159 VSS VSS nmos w=1u l=1u
M9665 n4156 n4022 net2910 VDD pmos w=2u l=1u
M9666 net2910 n4159 VDD VDD pmos w=2u l=1u
M9667 n4022 n4161 VSS VSS nmos w=1u l=1u
M9668 n4022 n4160 VSS VSS nmos w=1u l=1u
M9669 n4022 n4161 net2911 VDD pmos w=2u l=1u
M9670 net2911 n4160 VDD VDD pmos w=2u l=1u
M9671 n4159 net2912 VSS VSS nmos w=1u l=1u
M9672 net2913 n4160 VSS VSS nmos w=1u l=1u
M9673 net2912 n4161 net2913 VSS nmos w=1u l=1u
M9674 net2912 n4160 VDD VDD pmos w=2u l=1u
M9675 net2912 n4161 VDD VDD pmos w=2u l=1u
M9676 n4159 net2912 VDD VDD pmos w=2u l=1u
M9677 n4160 n4162 net2914 VSS nmos w=1u l=1u
M9678 net2914 n4044 VSS VSS nmos w=1u l=1u
M9679 n4160 n4162 VDD VDD pmos w=2u l=1u
M9680 n4160 n4044 VDD VDD pmos w=2u l=1u
M9681 n4162 N171 net2915 VSS nmos w=1u l=1u
M9682 net2915 n4163 VSS VSS nmos w=1u l=1u
M9683 n4162 N171 VDD VDD pmos w=2u l=1u
M9684 n4162 n4163 VDD VDD pmos w=2u l=1u
M9685 n4163 n3411 VSS VSS nmos w=1u l=1u
M9686 n4163 n4164 VSS VSS nmos w=1u l=1u
M9687 n4163 n3411 net2916 VDD pmos w=2u l=1u
M9688 net2916 n4164 VDD VDD pmos w=2u l=1u
M9689 n4044 n4165 net2917 VSS nmos w=1u l=1u
M9690 net2917 n4164 VSS VSS nmos w=1u l=1u
M9691 n4044 n4165 VDD VDD pmos w=2u l=1u
M9692 n4044 n4164 VDD VDD pmos w=2u l=1u
M9693 n4165 N307 net2918 VSS nmos w=1u l=1u
M9694 net2918 N171 VSS VSS nmos w=1u l=1u
M9695 n4165 N307 VDD VDD pmos w=2u l=1u
M9696 n4165 N171 VDD VDD pmos w=2u l=1u
M9697 n4164 net2919 VSS VSS nmos w=1u l=1u
M9698 net2920 n4166 VSS VSS nmos w=1u l=1u
M9699 net2919 n4045 net2920 VSS nmos w=1u l=1u
M9700 net2919 n4166 VDD VDD pmos w=2u l=1u
M9701 net2919 n4045 VDD VDD pmos w=2u l=1u
M9702 n4164 net2919 VDD VDD pmos w=2u l=1u
M9703 n4166 net2921 VSS VSS nmos w=1u l=1u
M9704 net2921 n4167 VSS VSS nmos w=1u l=1u
M9705 net2921 n4037 VSS VSS nmos w=1u l=1u
M9706 net2921 n4037 net2922 VDD pmos w=2u l=1u
M9707 n4166 net2921 VDD VDD pmos w=2u l=1u
M9708 net2922 n4167 VDD VDD pmos w=2u l=1u
M9709 n4037 n4038 VDD VDD pmos w=2u l=1u
M9710 n4037 n4038 VSS VSS nmos w=1u l=1u
M9711 n4045 n4168 net2923 VSS nmos w=1u l=1u
M9712 net2923 n4167 VSS VSS nmos w=1u l=1u
M9713 n4045 n4168 VDD VDD pmos w=2u l=1u
M9714 n4045 n4167 VDD VDD pmos w=2u l=1u
M9715 n4168 n4038 net2924 VSS nmos w=1u l=1u
M9716 net2924 n4169 VSS VSS nmos w=1u l=1u
M9717 n4168 n4038 VDD VDD pmos w=2u l=1u
M9718 n4168 n4169 VDD VDD pmos w=2u l=1u
M9719 n4038 N205 net2925 VSS nmos w=1u l=1u
M9720 net2925 n4170 VSS VSS nmos w=1u l=1u
M9721 n4038 N205 VDD VDD pmos w=2u l=1u
M9722 n4038 n4170 VDD VDD pmos w=2u l=1u
M9723 n4170 net2926 VSS VSS nmos w=1u l=1u
M9724 net2927 N188 VSS VSS nmos w=1u l=1u
M9725 net2926 n3741 net2927 VSS nmos w=1u l=1u
M9726 net2926 N188 VDD VDD pmos w=2u l=1u
M9727 net2926 n3741 VDD VDD pmos w=2u l=1u
M9728 n4170 net2926 VDD VDD pmos w=2u l=1u
M9729 n4169 n4172 net2928 VSS nmos w=1u l=1u
M9730 net2928 n4171 VSS VSS nmos w=1u l=1u
M9731 n4169 n4172 VDD VDD pmos w=2u l=1u
M9732 n4169 n4171 VDD VDD pmos w=2u l=1u
M9733 n4172 N273 net2929 VSS nmos w=1u l=1u
M9734 net2929 N205 VSS VSS nmos w=1u l=1u
M9735 n4172 N273 VDD VDD pmos w=2u l=1u
M9736 n4172 N205 VDD VDD pmos w=2u l=1u
M9737 n4171 N290 net2930 VSS nmos w=1u l=1u
M9738 net2930 N188 VSS VSS nmos w=1u l=1u
M9739 n4171 N290 VDD VDD pmos w=2u l=1u
M9740 n4171 N188 VDD VDD pmos w=2u l=1u
M9741 n4161 net2931 VSS VSS nmos w=1u l=1u
M9742 net2932 n4174 VSS VSS nmos w=1u l=1u
M9743 net2931 n4173 net2932 VSS nmos w=1u l=1u
M9744 net2931 n4174 VDD VDD pmos w=2u l=1u
M9745 net2931 n4173 VDD VDD pmos w=2u l=1u
M9746 n4161 net2931 VDD VDD pmos w=2u l=1u
M9747 n4154 n4151 VSS VSS nmos w=1u l=1u
M9748 n4154 n4152 VSS VSS nmos w=1u l=1u
M9749 n4154 n4151 net2933 VDD pmos w=2u l=1u
M9750 net2933 n4152 VDD VDD pmos w=2u l=1u
M9751 n4151 n4175 VDD VDD pmos w=2u l=1u
M9752 n4151 n4175 VSS VSS nmos w=1u l=1u
M9753 n4146 n4177 VSS VSS nmos w=1u l=1u
M9754 n4146 n4176 VSS VSS nmos w=1u l=1u
M9755 n4146 n4177 net2934 VDD pmos w=2u l=1u
M9756 net2934 n4176 VDD VDD pmos w=2u l=1u
M9757 n4177 net2935 VSS VSS nmos w=1u l=1u
M9758 net2936 n4143 VSS VSS nmos w=1u l=1u
M9759 net2935 n4144 net2936 VSS nmos w=1u l=1u
M9760 net2935 n4143 VDD VDD pmos w=2u l=1u
M9761 net2935 n4144 VDD VDD pmos w=2u l=1u
M9762 n4177 net2935 VDD VDD pmos w=2u l=1u
M9763 n4176 n4142 VDD VDD pmos w=2u l=1u
M9764 n4176 n4142 VSS VSS nmos w=1u l=1u
M9765 n4136 n4179 VSS VSS nmos w=1u l=1u
M9766 n4136 n4178 VSS VSS nmos w=1u l=1u
M9767 n4136 n4179 net2937 VDD pmos w=2u l=1u
M9768 net2937 n4178 VDD VDD pmos w=2u l=1u
M9769 n4179 n4133 VSS VSS nmos w=1u l=1u
M9770 n4179 n4134 VSS VSS nmos w=1u l=1u
M9771 n4179 n4133 net2938 VDD pmos w=2u l=1u
M9772 net2938 n4134 VDD VDD pmos w=2u l=1u
M9773 n4178 n4132 VDD VDD pmos w=2u l=1u
M9774 n4178 n4132 VSS VSS nmos w=1u l=1u
M9775 n4126 n4181 VSS VSS nmos w=1u l=1u
M9776 n4126 n4180 VSS VSS nmos w=1u l=1u
M9777 n4126 n4181 net2939 VDD pmos w=2u l=1u
M9778 net2939 n4180 VDD VDD pmos w=2u l=1u
M9779 n4181 net2940 VSS VSS nmos w=1u l=1u
M9780 net2941 n4123 VSS VSS nmos w=1u l=1u
M9781 net2940 n4124 net2941 VSS nmos w=1u l=1u
M9782 net2940 n4123 VDD VDD pmos w=2u l=1u
M9783 net2940 n4124 VDD VDD pmos w=2u l=1u
M9784 n4181 net2940 VDD VDD pmos w=2u l=1u
M9785 n4180 n4122 VDD VDD pmos w=2u l=1u
M9786 n4180 n4122 VSS VSS nmos w=1u l=1u
M9787 n4116 n4183 VSS VSS nmos w=1u l=1u
M9788 n4116 n4182 VSS VSS nmos w=1u l=1u
M9789 n4116 n4183 net2942 VDD pmos w=2u l=1u
M9790 net2942 n4182 VDD VDD pmos w=2u l=1u
M9791 n4183 net2943 VSS VSS nmos w=1u l=1u
M9792 net2944 n4113 VSS VSS nmos w=1u l=1u
M9793 net2943 n4114 net2944 VSS nmos w=1u l=1u
M9794 net2943 n4113 VDD VDD pmos w=2u l=1u
M9795 net2943 n4114 VDD VDD pmos w=2u l=1u
M9796 n4183 net2943 VDD VDD pmos w=2u l=1u
M9797 n4182 n4112 VDD VDD pmos w=2u l=1u
M9798 n4182 n4112 VSS VSS nmos w=1u l=1u
M9799 n4106 n4185 VSS VSS nmos w=1u l=1u
M9800 n4106 n4184 VSS VSS nmos w=1u l=1u
M9801 n4106 n4185 net2945 VDD pmos w=2u l=1u
M9802 net2945 n4184 VDD VDD pmos w=2u l=1u
M9803 n4185 net2946 VSS VSS nmos w=1u l=1u
M9804 net2947 n4103 VSS VSS nmos w=1u l=1u
M9805 net2946 n4104 net2947 VSS nmos w=1u l=1u
M9806 net2946 n4103 VDD VDD pmos w=2u l=1u
M9807 net2946 n4104 VDD VDD pmos w=2u l=1u
M9808 n4185 net2946 VDD VDD pmos w=2u l=1u
M9809 n4184 n4102 VDD VDD pmos w=2u l=1u
M9810 n4184 n4102 VSS VSS nmos w=1u l=1u
M9811 n4096 n4187 VSS VSS nmos w=1u l=1u
M9812 n4096 n4186 VSS VSS nmos w=1u l=1u
M9813 n4096 n4187 net2948 VDD pmos w=2u l=1u
M9814 net2948 n4186 VDD VDD pmos w=2u l=1u
M9815 n4187 n4189 VSS VSS nmos w=1u l=1u
M9816 n4187 n4188 VSS VSS nmos w=1u l=1u
M9817 n4187 n4189 net2949 VDD pmos w=2u l=1u
M9818 net2949 n4188 VDD VDD pmos w=2u l=1u
M9819 n4188 n4094 VDD VDD pmos w=2u l=1u
M9820 n4188 n4094 VSS VSS nmos w=1u l=1u
M9821 n4186 n4092 VDD VDD pmos w=2u l=1u
M9822 n4186 n4092 VSS VSS nmos w=1u l=1u
M9823 n4086 n4191 VSS VSS nmos w=1u l=1u
M9824 n4086 n4190 VSS VSS nmos w=1u l=1u
M9825 n4086 n4191 net2950 VDD pmos w=2u l=1u
M9826 net2950 n4190 VDD VDD pmos w=2u l=1u
M9827 n4191 n4193 VSS VSS nmos w=1u l=1u
M9828 n4191 n4192 VSS VSS nmos w=1u l=1u
M9829 n4191 n4193 net2951 VDD pmos w=2u l=1u
M9830 net2951 n4192 VDD VDD pmos w=2u l=1u
M9831 n4192 n4085 VDD VDD pmos w=2u l=1u
M9832 n4192 n4085 VSS VSS nmos w=1u l=1u
M9833 n4190 n4083 VDD VDD pmos w=2u l=1u
M9834 n4190 n4083 VSS VSS nmos w=1u l=1u
M9835 n4077 n4195 VSS VSS nmos w=1u l=1u
M9836 n4077 n4194 VSS VSS nmos w=1u l=1u
M9837 n4077 n4195 net2952 VDD pmos w=2u l=1u
M9838 net2952 n4194 VDD VDD pmos w=2u l=1u
M9839 n4195 n4075 VSS VSS nmos w=1u l=1u
M9840 n4195 n4076 VSS VSS nmos w=1u l=1u
M9841 n4195 n4075 net2953 VDD pmos w=2u l=1u
M9842 net2953 n4076 VDD VDD pmos w=2u l=1u
M9843 n4194 n4074 VDD VDD pmos w=2u l=1u
M9844 n4194 n4074 VSS VSS nmos w=1u l=1u
M9845 net2954 n4076 VSS VSS nmos w=1u l=1u
M9846 net2955 n4196 VSS VSS nmos w=1u l=1u
M9847 N4946 net2956 VSS VSS nmos w=1u l=1u
M9848 net2956 n4076 net2957 VSS nmos w=1u l=1u
M9849 net2956 net2954 net2955 VSS nmos w=1u l=1u
M9850 net2957 net2955 VSS VSS nmos w=1u l=1u
M9851 net2956 net2954 net2958 VDD pmos w=2u l=1u
M9852 net2954 n4076 VDD VDD pmos w=2u l=1u
M9853 net2955 n4076 net2956 VDD pmos w=2u l=1u
M9854 net2955 n4196 VDD VDD pmos w=2u l=1u
M9855 N4946 net2956 VDD VDD pmos w=2u l=1u
M9856 net2958 net2955 VDD VDD pmos w=2u l=1u
M9857 n4076 n2377 VSS VSS nmos w=1u l=1u
M9858 n4076 n3929 VSS VSS nmos w=1u l=1u
M9859 n4076 n2377 net2959 VDD pmos w=2u l=1u
M9860 net2959 n3929 VDD VDD pmos w=2u l=1u
M9861 n2377 N460 VDD VDD pmos w=2u l=1u
M9862 n2377 N460 VSS VSS nmos w=1u l=1u
M9863 n4196 n4075 VDD VDD pmos w=2u l=1u
M9864 n4196 n4075 VSS VSS nmos w=1u l=1u
M9865 n4075 n4074 net2960 VSS nmos w=1u l=1u
M9866 net2960 n4197 VSS VSS nmos w=1u l=1u
M9867 n4075 n4074 VDD VDD pmos w=2u l=1u
M9868 n4075 n4197 VDD VDD pmos w=2u l=1u
M9869 n4074 n4199 net2961 VSS nmos w=1u l=1u
M9870 net2961 n4198 VSS VSS nmos w=1u l=1u
M9871 n4074 n4199 VDD VDD pmos w=2u l=1u
M9872 n4074 n4198 VDD VDD pmos w=2u l=1u
M9873 n4199 n4201 net2962 VSS nmos w=1u l=1u
M9874 net2962 n4200 VSS VSS nmos w=1u l=1u
M9875 n4199 n4201 VDD VDD pmos w=2u l=1u
M9876 n4199 n4200 VDD VDD pmos w=2u l=1u
M9877 n4200 net2963 VSS VSS nmos w=1u l=1u
M9878 net2963 n4202 VSS VSS nmos w=1u l=1u
M9879 net2963 n4203 VSS VSS nmos w=1u l=1u
M9880 net2963 n4203 net2964 VDD pmos w=2u l=1u
M9881 n4200 net2963 VDD VDD pmos w=2u l=1u
M9882 net2964 n4202 VDD VDD pmos w=2u l=1u
M9883 net2965 n4084 VSS VSS nmos w=1u l=1u
M9884 net2966 n4085 VSS VSS nmos w=1u l=1u
M9885 n4198 net2967 VSS VSS nmos w=1u l=1u
M9886 net2967 n4084 net2968 VSS nmos w=1u l=1u
M9887 net2967 net2965 net2966 VSS nmos w=1u l=1u
M9888 net2968 net2966 VSS VSS nmos w=1u l=1u
M9889 net2967 net2965 net2969 VDD pmos w=2u l=1u
M9890 net2965 n4084 VDD VDD pmos w=2u l=1u
M9891 net2966 n4084 net2967 VDD pmos w=2u l=1u
M9892 net2966 n4085 VDD VDD pmos w=2u l=1u
M9893 n4198 net2967 VDD VDD pmos w=2u l=1u
M9894 net2969 net2966 VDD VDD pmos w=2u l=1u
M9895 n4084 n4193 VDD VDD pmos w=2u l=1u
M9896 n4084 n4193 VSS VSS nmos w=1u l=1u
M9897 n4197 n4205 net2970 VSS nmos w=1u l=1u
M9898 net2970 n4204 VSS VSS nmos w=1u l=1u
M9899 n4197 n4205 VDD VDD pmos w=2u l=1u
M9900 n4197 n4204 VDD VDD pmos w=2u l=1u
M9901 net2971 n4085 VSS VSS nmos w=1u l=1u
M9902 net2972 n4193 VSS VSS nmos w=1u l=1u
M9903 n4205 net2973 VSS VSS nmos w=1u l=1u
M9904 net2973 n4085 net2974 VSS nmos w=1u l=1u
M9905 net2973 net2971 net2972 VSS nmos w=1u l=1u
M9906 net2974 net2972 VSS VSS nmos w=1u l=1u
M9907 net2973 net2971 net2975 VDD pmos w=2u l=1u
M9908 net2971 n4085 VDD VDD pmos w=2u l=1u
M9909 net2972 n4085 net2973 VDD pmos w=2u l=1u
M9910 net2972 n4193 VDD VDD pmos w=2u l=1u
M9911 n4205 net2973 VDD VDD pmos w=2u l=1u
M9912 net2975 net2972 VDD VDD pmos w=2u l=1u
M9913 n4085 N443 net2976 VSS nmos w=1u l=1u
M9914 net2976 N18 VSS VSS nmos w=1u l=1u
M9915 n4085 N443 VDD VDD pmos w=2u l=1u
M9916 n4085 N18 VDD VDD pmos w=2u l=1u
M9917 n4193 n4083 net2977 VSS nmos w=1u l=1u
M9918 net2977 n4206 VSS VSS nmos w=1u l=1u
M9919 n4193 n4083 VDD VDD pmos w=2u l=1u
M9920 n4193 n4206 VDD VDD pmos w=2u l=1u
M9921 n4083 n4208 net2978 VSS nmos w=1u l=1u
M9922 net2978 n4207 VSS VSS nmos w=1u l=1u
M9923 n4083 n4208 VDD VDD pmos w=2u l=1u
M9924 n4083 n4207 VDD VDD pmos w=2u l=1u
M9925 n4208 n4210 net2979 VSS nmos w=1u l=1u
M9926 net2979 n4209 VSS VSS nmos w=1u l=1u
M9927 n4208 n4210 VDD VDD pmos w=2u l=1u
M9928 n4208 n4209 VDD VDD pmos w=2u l=1u
M9929 n4209 n4212 net2980 VSS nmos w=1u l=1u
M9930 net2980 n4211 VSS VSS nmos w=1u l=1u
M9931 n4209 n4212 VDD VDD pmos w=2u l=1u
M9932 n4209 n4211 VDD VDD pmos w=2u l=1u
M9933 net2981 n4093 VSS VSS nmos w=1u l=1u
M9934 net2982 n4094 VSS VSS nmos w=1u l=1u
M9935 n4207 net2983 VSS VSS nmos w=1u l=1u
M9936 net2983 n4093 net2984 VSS nmos w=1u l=1u
M9937 net2983 net2981 net2982 VSS nmos w=1u l=1u
M9938 net2984 net2982 VSS VSS nmos w=1u l=1u
M9939 net2983 net2981 net2985 VDD pmos w=2u l=1u
M9940 net2981 n4093 VDD VDD pmos w=2u l=1u
M9941 net2982 n4093 net2983 VDD pmos w=2u l=1u
M9942 net2982 n4094 VDD VDD pmos w=2u l=1u
M9943 n4207 net2983 VDD VDD pmos w=2u l=1u
M9944 net2985 net2982 VDD VDD pmos w=2u l=1u
M9945 n4093 n4189 VDD VDD pmos w=2u l=1u
M9946 n4093 n4189 VSS VSS nmos w=1u l=1u
M9947 n4206 n4214 net2986 VSS nmos w=1u l=1u
M9948 net2986 n4213 VSS VSS nmos w=1u l=1u
M9949 n4206 n4214 VDD VDD pmos w=2u l=1u
M9950 n4206 n4213 VDD VDD pmos w=2u l=1u
M9951 net2987 n4094 VSS VSS nmos w=1u l=1u
M9952 net2988 n4189 VSS VSS nmos w=1u l=1u
M9953 n4214 net2989 VSS VSS nmos w=1u l=1u
M9954 net2989 n4094 net2990 VSS nmos w=1u l=1u
M9955 net2989 net2987 net2988 VSS nmos w=1u l=1u
M9956 net2990 net2988 VSS VSS nmos w=1u l=1u
M9957 net2989 net2987 net2991 VDD pmos w=2u l=1u
M9958 net2987 n4094 VDD VDD pmos w=2u l=1u
M9959 net2988 n4094 net2989 VDD pmos w=2u l=1u
M9960 net2988 n4189 VDD VDD pmos w=2u l=1u
M9961 n4214 net2989 VDD VDD pmos w=2u l=1u
M9962 net2991 net2988 VDD VDD pmos w=2u l=1u
M9963 n4094 N426 net2992 VSS nmos w=1u l=1u
M9964 net2992 N35 VSS VSS nmos w=1u l=1u
M9965 n4094 N426 VDD VDD pmos w=2u l=1u
M9966 n4094 N35 VDD VDD pmos w=2u l=1u
M9967 n4189 n4092 net2993 VSS nmos w=1u l=1u
M9968 net2993 n4215 VSS VSS nmos w=1u l=1u
M9969 n4189 n4092 VDD VDD pmos w=2u l=1u
M9970 n4189 n4215 VDD VDD pmos w=2u l=1u
M9971 n4092 n4217 net2994 VSS nmos w=1u l=1u
M9972 net2994 n4216 VSS VSS nmos w=1u l=1u
M9973 n4092 n4217 VDD VDD pmos w=2u l=1u
M9974 n4092 n4216 VDD VDD pmos w=2u l=1u
M9975 n4217 n4219 net2995 VSS nmos w=1u l=1u
M9976 net2995 n4218 VSS VSS nmos w=1u l=1u
M9977 n4217 n4219 VDD VDD pmos w=2u l=1u
M9978 n4217 n4218 VDD VDD pmos w=2u l=1u
M9979 n4218 n4221 net2996 VSS nmos w=1u l=1u
M9980 net2996 n4220 VSS VSS nmos w=1u l=1u
M9981 n4218 n4221 VDD VDD pmos w=2u l=1u
M9982 n4218 n4220 VDD VDD pmos w=2u l=1u
M9983 net2997 n4103 VSS VSS nmos w=1u l=1u
M9984 net2998 n4104 VSS VSS nmos w=1u l=1u
M9985 n4216 net2999 VSS VSS nmos w=1u l=1u
M9986 net2999 n4103 net3000 VSS nmos w=1u l=1u
M9987 net2999 net2997 net2998 VSS nmos w=1u l=1u
M9988 net3000 net2998 VSS VSS nmos w=1u l=1u
M9989 net2999 net2997 net3001 VDD pmos w=2u l=1u
M9990 net2997 n4103 VDD VDD pmos w=2u l=1u
M9991 net2998 n4103 net2999 VDD pmos w=2u l=1u
M9992 net2998 n4104 VDD VDD pmos w=2u l=1u
M9993 n4216 net2999 VDD VDD pmos w=2u l=1u
M9994 net3001 net2998 VDD VDD pmos w=2u l=1u
M9995 n4103 n4222 VDD VDD pmos w=2u l=1u
M9996 n4103 n4222 VSS VSS nmos w=1u l=1u
M9997 n4215 n4224 net3002 VSS nmos w=1u l=1u
M9998 net3002 n4223 VSS VSS nmos w=1u l=1u
M9999 n4215 n4224 VDD VDD pmos w=2u l=1u
M10000 n4215 n4223 VDD VDD pmos w=2u l=1u
M10001 net3003 n4104 VSS VSS nmos w=1u l=1u
M10002 net3004 n4222 VSS VSS nmos w=1u l=1u
M10003 n4224 net3005 VSS VSS nmos w=1u l=1u
M10004 net3005 n4104 net3006 VSS nmos w=1u l=1u
M10005 net3005 net3003 net3004 VSS nmos w=1u l=1u
M10006 net3006 net3004 VSS VSS nmos w=1u l=1u
M10007 net3005 net3003 net3007 VDD pmos w=2u l=1u
M10008 net3003 n4104 VDD VDD pmos w=2u l=1u
M10009 net3004 n4104 net3005 VDD pmos w=2u l=1u
M10010 net3004 n4222 VDD VDD pmos w=2u l=1u
M10011 n4224 net3005 VDD VDD pmos w=2u l=1u
M10012 net3007 net3004 VDD VDD pmos w=2u l=1u
M10013 n4104 N409 net3008 VSS nmos w=1u l=1u
M10014 net3008 N52 VSS VSS nmos w=1u l=1u
M10015 n4104 N409 VDD VDD pmos w=2u l=1u
M10016 n4104 N52 VDD VDD pmos w=2u l=1u
M10017 n4222 n4102 net3009 VSS nmos w=1u l=1u
M10018 net3009 n4225 VSS VSS nmos w=1u l=1u
M10019 n4222 n4102 VDD VDD pmos w=2u l=1u
M10020 n4222 n4225 VDD VDD pmos w=2u l=1u
M10021 n4102 n4227 net3010 VSS nmos w=1u l=1u
M10022 net3010 n4226 VSS VSS nmos w=1u l=1u
M10023 n4102 n4227 VDD VDD pmos w=2u l=1u
M10024 n4102 n4226 VDD VDD pmos w=2u l=1u
M10025 n4227 n4229 net3011 VSS nmos w=1u l=1u
M10026 net3011 n4228 VSS VSS nmos w=1u l=1u
M10027 n4227 n4229 VDD VDD pmos w=2u l=1u
M10028 n4227 n4228 VDD VDD pmos w=2u l=1u
M10029 n4228 n4231 net3012 VSS nmos w=1u l=1u
M10030 net3012 n4230 VSS VSS nmos w=1u l=1u
M10031 n4228 n4231 VDD VDD pmos w=2u l=1u
M10032 n4228 n4230 VDD VDD pmos w=2u l=1u
M10033 net3013 n4113 VSS VSS nmos w=1u l=1u
M10034 net3014 n4114 VSS VSS nmos w=1u l=1u
M10035 n4226 net3015 VSS VSS nmos w=1u l=1u
M10036 net3015 n4113 net3016 VSS nmos w=1u l=1u
M10037 net3015 net3013 net3014 VSS nmos w=1u l=1u
M10038 net3016 net3014 VSS VSS nmos w=1u l=1u
M10039 net3015 net3013 net3017 VDD pmos w=2u l=1u
M10040 net3013 n4113 VDD VDD pmos w=2u l=1u
M10041 net3014 n4113 net3015 VDD pmos w=2u l=1u
M10042 net3014 n4114 VDD VDD pmos w=2u l=1u
M10043 n4226 net3015 VDD VDD pmos w=2u l=1u
M10044 net3017 net3014 VDD VDD pmos w=2u l=1u
M10045 n4113 n4232 VDD VDD pmos w=2u l=1u
M10046 n4113 n4232 VSS VSS nmos w=1u l=1u
M10047 n4225 n4234 net3018 VSS nmos w=1u l=1u
M10048 net3018 n4233 VSS VSS nmos w=1u l=1u
M10049 n4225 n4234 VDD VDD pmos w=2u l=1u
M10050 n4225 n4233 VDD VDD pmos w=2u l=1u
M10051 net3019 n4114 VSS VSS nmos w=1u l=1u
M10052 net3020 n4232 VSS VSS nmos w=1u l=1u
M10053 n4234 net3021 VSS VSS nmos w=1u l=1u
M10054 net3021 n4114 net3022 VSS nmos w=1u l=1u
M10055 net3021 net3019 net3020 VSS nmos w=1u l=1u
M10056 net3022 net3020 VSS VSS nmos w=1u l=1u
M10057 net3021 net3019 net3023 VDD pmos w=2u l=1u
M10058 net3019 n4114 VDD VDD pmos w=2u l=1u
M10059 net3020 n4114 net3021 VDD pmos w=2u l=1u
M10060 net3020 n4232 VDD VDD pmos w=2u l=1u
M10061 n4234 net3021 VDD VDD pmos w=2u l=1u
M10062 net3023 net3020 VDD VDD pmos w=2u l=1u
M10063 n4114 N392 net3024 VSS nmos w=1u l=1u
M10064 net3024 N69 VSS VSS nmos w=1u l=1u
M10065 n4114 N392 VDD VDD pmos w=2u l=1u
M10066 n4114 N69 VDD VDD pmos w=2u l=1u
M10067 n4232 n4112 net3025 VSS nmos w=1u l=1u
M10068 net3025 n4235 VSS VSS nmos w=1u l=1u
M10069 n4232 n4112 VDD VDD pmos w=2u l=1u
M10070 n4232 n4235 VDD VDD pmos w=2u l=1u
M10071 n4112 n4237 net3026 VSS nmos w=1u l=1u
M10072 net3026 n4236 VSS VSS nmos w=1u l=1u
M10073 n4112 n4237 VDD VDD pmos w=2u l=1u
M10074 n4112 n4236 VDD VDD pmos w=2u l=1u
M10075 n4237 n4239 net3027 VSS nmos w=1u l=1u
M10076 net3027 n4238 VSS VSS nmos w=1u l=1u
M10077 n4237 n4239 VDD VDD pmos w=2u l=1u
M10078 n4237 n4238 VDD VDD pmos w=2u l=1u
M10079 n4238 n4241 net3028 VSS nmos w=1u l=1u
M10080 net3028 n4240 VSS VSS nmos w=1u l=1u
M10081 n4238 n4241 VDD VDD pmos w=2u l=1u
M10082 n4238 n4240 VDD VDD pmos w=2u l=1u
M10083 net3029 n4123 VSS VSS nmos w=1u l=1u
M10084 net3030 n4124 VSS VSS nmos w=1u l=1u
M10085 n4236 net3031 VSS VSS nmos w=1u l=1u
M10086 net3031 n4123 net3032 VSS nmos w=1u l=1u
M10087 net3031 net3029 net3030 VSS nmos w=1u l=1u
M10088 net3032 net3030 VSS VSS nmos w=1u l=1u
M10089 net3031 net3029 net3033 VDD pmos w=2u l=1u
M10090 net3029 n4123 VDD VDD pmos w=2u l=1u
M10091 net3030 n4123 net3031 VDD pmos w=2u l=1u
M10092 net3030 n4124 VDD VDD pmos w=2u l=1u
M10093 n4236 net3031 VDD VDD pmos w=2u l=1u
M10094 net3033 net3030 VDD VDD pmos w=2u l=1u
M10095 n4123 n4242 VDD VDD pmos w=2u l=1u
M10096 n4123 n4242 VSS VSS nmos w=1u l=1u
M10097 n4235 n4244 net3034 VSS nmos w=1u l=1u
M10098 net3034 n4243 VSS VSS nmos w=1u l=1u
M10099 n4235 n4244 VDD VDD pmos w=2u l=1u
M10100 n4235 n4243 VDD VDD pmos w=2u l=1u
M10101 net3035 n4124 VSS VSS nmos w=1u l=1u
M10102 net3036 n4242 VSS VSS nmos w=1u l=1u
M10103 n4244 net3037 VSS VSS nmos w=1u l=1u
M10104 net3037 n4124 net3038 VSS nmos w=1u l=1u
M10105 net3037 net3035 net3036 VSS nmos w=1u l=1u
M10106 net3038 net3036 VSS VSS nmos w=1u l=1u
M10107 net3037 net3035 net3039 VDD pmos w=2u l=1u
M10108 net3035 n4124 VDD VDD pmos w=2u l=1u
M10109 net3036 n4124 net3037 VDD pmos w=2u l=1u
M10110 net3036 n4242 VDD VDD pmos w=2u l=1u
M10111 n4244 net3037 VDD VDD pmos w=2u l=1u
M10112 net3039 net3036 VDD VDD pmos w=2u l=1u
M10113 n4124 N375 net3040 VSS nmos w=1u l=1u
M10114 net3040 N86 VSS VSS nmos w=1u l=1u
M10115 n4124 N375 VDD VDD pmos w=2u l=1u
M10116 n4124 N86 VDD VDD pmos w=2u l=1u
M10117 n4242 n4122 net3041 VSS nmos w=1u l=1u
M10118 net3041 n4245 VSS VSS nmos w=1u l=1u
M10119 n4242 n4122 VDD VDD pmos w=2u l=1u
M10120 n4242 n4245 VDD VDD pmos w=2u l=1u
M10121 n4122 n4247 net3042 VSS nmos w=1u l=1u
M10122 net3042 n4246 VSS VSS nmos w=1u l=1u
M10123 n4122 n4247 VDD VDD pmos w=2u l=1u
M10124 n4122 n4246 VDD VDD pmos w=2u l=1u
M10125 n4247 n4249 net3043 VSS nmos w=1u l=1u
M10126 net3043 n4248 VSS VSS nmos w=1u l=1u
M10127 n4247 n4249 VDD VDD pmos w=2u l=1u
M10128 n4247 n4248 VDD VDD pmos w=2u l=1u
M10129 n4248 net3044 VSS VSS nmos w=1u l=1u
M10130 net3044 n4250 VSS VSS nmos w=1u l=1u
M10131 net3044 n4251 VSS VSS nmos w=1u l=1u
M10132 net3044 n4251 net3045 VDD pmos w=2u l=1u
M10133 n4248 net3044 VDD VDD pmos w=2u l=1u
M10134 net3045 n4250 VDD VDD pmos w=2u l=1u
M10135 net3046 n4133 VSS VSS nmos w=1u l=1u
M10136 net3047 n4134 VSS VSS nmos w=1u l=1u
M10137 n4246 net3048 VSS VSS nmos w=1u l=1u
M10138 net3048 n4133 net3049 VSS nmos w=1u l=1u
M10139 net3048 net3046 net3047 VSS nmos w=1u l=1u
M10140 net3049 net3047 VSS VSS nmos w=1u l=1u
M10141 net3048 net3046 net3050 VDD pmos w=2u l=1u
M10142 net3046 n4133 VDD VDD pmos w=2u l=1u
M10143 net3047 n4133 net3048 VDD pmos w=2u l=1u
M10144 net3047 n4134 VDD VDD pmos w=2u l=1u
M10145 n4246 net3048 VDD VDD pmos w=2u l=1u
M10146 net3050 net3047 VDD VDD pmos w=2u l=1u
M10147 n4134 n4252 VDD VDD pmos w=2u l=1u
M10148 n4134 n4252 VSS VSS nmos w=1u l=1u
M10149 n4245 n4254 net3051 VSS nmos w=1u l=1u
M10150 net3051 n4253 VSS VSS nmos w=1u l=1u
M10151 n4245 n4254 VDD VDD pmos w=2u l=1u
M10152 n4245 n4253 VDD VDD pmos w=2u l=1u
M10153 net3052 n4252 VSS VSS nmos w=1u l=1u
M10154 net3053 n4133 VSS VSS nmos w=1u l=1u
M10155 n4254 net3054 VSS VSS nmos w=1u l=1u
M10156 net3054 n4252 net3055 VSS nmos w=1u l=1u
M10157 net3054 net3052 net3053 VSS nmos w=1u l=1u
M10158 net3055 net3053 VSS VSS nmos w=1u l=1u
M10159 net3054 net3052 net3056 VDD pmos w=2u l=1u
M10160 net3052 n4252 VDD VDD pmos w=2u l=1u
M10161 net3053 n4252 net3054 VDD pmos w=2u l=1u
M10162 net3053 n4133 VDD VDD pmos w=2u l=1u
M10163 n4254 net3054 VDD VDD pmos w=2u l=1u
M10164 net3056 net3053 VDD VDD pmos w=2u l=1u
M10165 n4252 N358 net3057 VSS nmos w=1u l=1u
M10166 net3057 N103 VSS VSS nmos w=1u l=1u
M10167 n4252 N358 VDD VDD pmos w=2u l=1u
M10168 n4252 N103 VDD VDD pmos w=2u l=1u
M10169 n4133 n4132 net3058 VSS nmos w=1u l=1u
M10170 net3058 n4255 VSS VSS nmos w=1u l=1u
M10171 n4133 n4132 VDD VDD pmos w=2u l=1u
M10172 n4133 n4255 VDD VDD pmos w=2u l=1u
M10173 n4132 n4257 net3059 VSS nmos w=1u l=1u
M10174 net3059 n4256 VSS VSS nmos w=1u l=1u
M10175 n4132 n4257 VDD VDD pmos w=2u l=1u
M10176 n4132 n4256 VDD VDD pmos w=2u l=1u
M10177 n4257 n4259 net3060 VSS nmos w=1u l=1u
M10178 net3060 n4258 VSS VSS nmos w=1u l=1u
M10179 n4257 n4259 VDD VDD pmos w=2u l=1u
M10180 n4257 n4258 VDD VDD pmos w=2u l=1u
M10181 n4258 n4261 net3061 VSS nmos w=1u l=1u
M10182 net3061 n4260 VSS VSS nmos w=1u l=1u
M10183 n4258 n4261 VDD VDD pmos w=2u l=1u
M10184 n4258 n4260 VDD VDD pmos w=2u l=1u
M10185 net3062 n4143 VSS VSS nmos w=1u l=1u
M10186 net3063 n4144 VSS VSS nmos w=1u l=1u
M10187 n4256 net3064 VSS VSS nmos w=1u l=1u
M10188 net3064 n4143 net3065 VSS nmos w=1u l=1u
M10189 net3064 net3062 net3063 VSS nmos w=1u l=1u
M10190 net3065 net3063 VSS VSS nmos w=1u l=1u
M10191 net3064 net3062 net3066 VDD pmos w=2u l=1u
M10192 net3062 n4143 VDD VDD pmos w=2u l=1u
M10193 net3063 n4143 net3064 VDD pmos w=2u l=1u
M10194 net3063 n4144 VDD VDD pmos w=2u l=1u
M10195 n4256 net3064 VDD VDD pmos w=2u l=1u
M10196 net3066 net3063 VDD VDD pmos w=2u l=1u
M10197 n4143 n4262 VDD VDD pmos w=2u l=1u
M10198 n4143 n4262 VSS VSS nmos w=1u l=1u
M10199 n4255 n4264 net3067 VSS nmos w=1u l=1u
M10200 net3067 n4263 VSS VSS nmos w=1u l=1u
M10201 n4255 n4264 VDD VDD pmos w=2u l=1u
M10202 n4255 n4263 VDD VDD pmos w=2u l=1u
M10203 net3068 n4144 VSS VSS nmos w=1u l=1u
M10204 net3069 n4262 VSS VSS nmos w=1u l=1u
M10205 n4264 net3070 VSS VSS nmos w=1u l=1u
M10206 net3070 n4144 net3071 VSS nmos w=1u l=1u
M10207 net3070 net3068 net3069 VSS nmos w=1u l=1u
M10208 net3071 net3069 VSS VSS nmos w=1u l=1u
M10209 net3070 net3068 net3072 VDD pmos w=2u l=1u
M10210 net3068 n4144 VDD VDD pmos w=2u l=1u
M10211 net3069 n4144 net3070 VDD pmos w=2u l=1u
M10212 net3069 n4262 VDD VDD pmos w=2u l=1u
M10213 n4264 net3070 VDD VDD pmos w=2u l=1u
M10214 net3072 net3069 VDD VDD pmos w=2u l=1u
M10215 n4144 N341 net3073 VSS nmos w=1u l=1u
M10216 net3073 N120 VSS VSS nmos w=1u l=1u
M10217 n4144 N341 VDD VDD pmos w=2u l=1u
M10218 n4144 N120 VDD VDD pmos w=2u l=1u
M10219 n4262 n4142 net3074 VSS nmos w=1u l=1u
M10220 net3074 n4265 VSS VSS nmos w=1u l=1u
M10221 n4262 n4142 VDD VDD pmos w=2u l=1u
M10222 n4262 n4265 VDD VDD pmos w=2u l=1u
M10223 n4142 n4267 net3075 VSS nmos w=1u l=1u
M10224 net3075 n4266 VSS VSS nmos w=1u l=1u
M10225 n4142 n4267 VDD VDD pmos w=2u l=1u
M10226 n4142 n4266 VDD VDD pmos w=2u l=1u
M10227 n4267 net3076 VSS VSS nmos w=1u l=1u
M10228 net3076 n4268 VSS VSS nmos w=1u l=1u
M10229 net3076 n4269 VSS VSS nmos w=1u l=1u
M10230 net3076 n4269 net3077 VDD pmos w=2u l=1u
M10231 n4267 net3076 VDD VDD pmos w=2u l=1u
M10232 net3077 n4268 VDD VDD pmos w=2u l=1u
M10233 n4266 net3078 VSS VSS nmos w=1u l=1u
M10234 net3079 n4270 VSS VSS nmos w=1u l=1u
M10235 net3078 n4175 net3079 VSS nmos w=1u l=1u
M10236 net3078 n4270 VDD VDD pmos w=2u l=1u
M10237 net3078 n4175 VDD VDD pmos w=2u l=1u
M10238 n4266 net3078 VDD VDD pmos w=2u l=1u
M10239 n4265 n4272 net3080 VSS nmos w=1u l=1u
M10240 net3080 n4271 VSS VSS nmos w=1u l=1u
M10241 n4265 n4272 VDD VDD pmos w=2u l=1u
M10242 n4265 n4271 VDD VDD pmos w=2u l=1u
M10243 n4272 n4175 net3081 VSS nmos w=1u l=1u
M10244 net3081 n4270 VSS VSS nmos w=1u l=1u
M10245 n4272 n4175 VDD VDD pmos w=2u l=1u
M10246 n4272 n4270 VDD VDD pmos w=2u l=1u
M10247 n4175 n4274 net3082 VSS nmos w=1u l=1u
M10248 net3082 n4273 VSS VSS nmos w=1u l=1u
M10249 n4175 n4274 VDD VDD pmos w=2u l=1u
M10250 n4175 n4273 VDD VDD pmos w=2u l=1u
M10251 n4274 N324 net3083 VSS nmos w=1u l=1u
M10252 net3083 N137 VSS VSS nmos w=1u l=1u
M10253 n4274 N324 VDD VDD pmos w=2u l=1u
M10254 n4274 N137 VDD VDD pmos w=2u l=1u
M10255 n4270 N137 net3084 VSS nmos w=1u l=1u
M10256 net3084 n4275 VSS VSS nmos w=1u l=1u
M10257 n4270 N137 VDD VDD pmos w=2u l=1u
M10258 n4270 n4275 VDD VDD pmos w=2u l=1u
M10259 n4275 n3257 VSS VSS nmos w=1u l=1u
M10260 n4275 n4273 VSS VSS nmos w=1u l=1u
M10261 n4275 n3257 net3085 VDD pmos w=2u l=1u
M10262 net3085 n4273 VDD VDD pmos w=2u l=1u
M10263 n4273 n4152 VSS VSS nmos w=1u l=1u
M10264 n4273 n4276 VSS VSS nmos w=1u l=1u
M10265 n4273 n4152 net3086 VDD pmos w=2u l=1u
M10266 net3086 n4276 VDD VDD pmos w=2u l=1u
M10267 n4152 n4278 VSS VSS nmos w=1u l=1u
M10268 n4152 n4277 VSS VSS nmos w=1u l=1u
M10269 n4152 n4278 net3087 VDD pmos w=2u l=1u
M10270 net3087 n4277 VDD VDD pmos w=2u l=1u
M10271 n4276 net3088 VSS VSS nmos w=1u l=1u
M10272 net3089 n4277 VSS VSS nmos w=1u l=1u
M10273 net3088 n4278 net3089 VSS nmos w=1u l=1u
M10274 net3088 n4277 VDD VDD pmos w=2u l=1u
M10275 net3088 n4278 VDD VDD pmos w=2u l=1u
M10276 n4276 net3088 VDD VDD pmos w=2u l=1u
M10277 n4277 n4279 net3090 VSS nmos w=1u l=1u
M10278 net3090 n4173 VSS VSS nmos w=1u l=1u
M10279 n4277 n4279 VDD VDD pmos w=2u l=1u
M10280 n4277 n4173 VDD VDD pmos w=2u l=1u
M10281 n4279 N154 net3091 VSS nmos w=1u l=1u
M10282 net3091 n4280 VSS VSS nmos w=1u l=1u
M10283 n4279 N154 VDD VDD pmos w=2u l=1u
M10284 n4279 n4280 VDD VDD pmos w=2u l=1u
M10285 n4280 n3411 VSS VSS nmos w=1u l=1u
M10286 n4280 n4281 VSS VSS nmos w=1u l=1u
M10287 n4280 n3411 net3092 VDD pmos w=2u l=1u
M10288 net3092 n4281 VDD VDD pmos w=2u l=1u
M10289 n4173 n4282 net3093 VSS nmos w=1u l=1u
M10290 net3093 n4281 VSS VSS nmos w=1u l=1u
M10291 n4173 n4282 VDD VDD pmos w=2u l=1u
M10292 n4173 n4281 VDD VDD pmos w=2u l=1u
M10293 n4282 N307 net3094 VSS nmos w=1u l=1u
M10294 net3094 N154 VSS VSS nmos w=1u l=1u
M10295 n4282 N307 VDD VDD pmos w=2u l=1u
M10296 n4282 N154 VDD VDD pmos w=2u l=1u
M10297 n4281 net3095 VSS VSS nmos w=1u l=1u
M10298 net3096 n4283 VSS VSS nmos w=1u l=1u
M10299 net3095 n4174 net3096 VSS nmos w=1u l=1u
M10300 net3095 n4283 VDD VDD pmos w=2u l=1u
M10301 net3095 n4174 VDD VDD pmos w=2u l=1u
M10302 n4281 net3095 VDD VDD pmos w=2u l=1u
M10303 n4283 n4167 net3097 VSS nmos w=1u l=1u
M10304 net3097 n4284 VSS VSS nmos w=1u l=1u
M10305 n4283 n4167 VDD VDD pmos w=2u l=1u
M10306 n4283 n4284 VDD VDD pmos w=2u l=1u
M10307 n4174 n4286 net3098 VSS nmos w=1u l=1u
M10308 net3098 n4285 VSS VSS nmos w=1u l=1u
M10309 n4174 n4286 VDD VDD pmos w=2u l=1u
M10310 n4174 n4285 VDD VDD pmos w=2u l=1u
M10311 n4286 n4167 net3099 VSS nmos w=1u l=1u
M10312 net3099 n4287 VSS VSS nmos w=1u l=1u
M10313 n4286 n4167 VDD VDD pmos w=2u l=1u
M10314 n4286 n4287 VDD VDD pmos w=2u l=1u
M10315 n4167 N188 net3100 VSS nmos w=1u l=1u
M10316 net3100 n4288 VSS VSS nmos w=1u l=1u
M10317 n4167 N188 VDD VDD pmos w=2u l=1u
M10318 n4167 n4288 VDD VDD pmos w=2u l=1u
M10319 n4288 net3101 VSS VSS nmos w=1u l=1u
M10320 net3102 N171 VSS VSS nmos w=1u l=1u
M10321 net3101 n3741 net3102 VSS nmos w=1u l=1u
M10322 net3101 N171 VDD VDD pmos w=2u l=1u
M10323 net3101 n3741 VDD VDD pmos w=2u l=1u
M10324 n4288 net3101 VDD VDD pmos w=2u l=1u
M10325 n4287 n4290 net3103 VSS nmos w=1u l=1u
M10326 net3103 n4289 VSS VSS nmos w=1u l=1u
M10327 n4287 n4290 VDD VDD pmos w=2u l=1u
M10328 n4287 n4289 VDD VDD pmos w=2u l=1u
M10329 n4290 N273 net3104 VSS nmos w=1u l=1u
M10330 net3104 N188 VSS VSS nmos w=1u l=1u
M10331 n4290 N273 VDD VDD pmos w=2u l=1u
M10332 n4290 N188 VDD VDD pmos w=2u l=1u
M10333 n4289 N290 net3105 VSS nmos w=1u l=1u
M10334 net3105 N171 VSS VSS nmos w=1u l=1u
M10335 n4289 N290 VDD VDD pmos w=2u l=1u
M10336 n4289 N171 VDD VDD pmos w=2u l=1u
M10337 n4278 net3106 VSS VSS nmos w=1u l=1u
M10338 net3107 n4292 VSS VSS nmos w=1u l=1u
M10339 net3106 n4291 net3107 VSS nmos w=1u l=1u
M10340 net3106 n4292 VDD VDD pmos w=2u l=1u
M10341 net3106 n4291 VDD VDD pmos w=2u l=1u
M10342 n4278 net3106 VDD VDD pmos w=2u l=1u
M10343 n4271 n4268 VSS VSS nmos w=1u l=1u
M10344 n4271 n4269 VSS VSS nmos w=1u l=1u
M10345 n4271 n4268 net3108 VDD pmos w=2u l=1u
M10346 net3108 n4269 VDD VDD pmos w=2u l=1u
M10347 n4268 n4293 VDD VDD pmos w=2u l=1u
M10348 n4268 n4293 VSS VSS nmos w=1u l=1u
M10349 n4263 n4295 VSS VSS nmos w=1u l=1u
M10350 n4263 n4294 VSS VSS nmos w=1u l=1u
M10351 n4263 n4295 net3109 VDD pmos w=2u l=1u
M10352 net3109 n4294 VDD VDD pmos w=2u l=1u
M10353 n4295 net3110 VSS VSS nmos w=1u l=1u
M10354 net3111 n4260 VSS VSS nmos w=1u l=1u
M10355 net3110 n4261 net3111 VSS nmos w=1u l=1u
M10356 net3110 n4260 VDD VDD pmos w=2u l=1u
M10357 net3110 n4261 VDD VDD pmos w=2u l=1u
M10358 n4295 net3110 VDD VDD pmos w=2u l=1u
M10359 n4294 n4259 VDD VDD pmos w=2u l=1u
M10360 n4294 n4259 VSS VSS nmos w=1u l=1u
M10361 n4253 n4297 VSS VSS nmos w=1u l=1u
M10362 n4253 n4296 VSS VSS nmos w=1u l=1u
M10363 n4253 n4297 net3112 VDD pmos w=2u l=1u
M10364 net3112 n4296 VDD VDD pmos w=2u l=1u
M10365 n4297 n4250 VSS VSS nmos w=1u l=1u
M10366 n4297 n4251 VSS VSS nmos w=1u l=1u
M10367 n4297 n4250 net3113 VDD pmos w=2u l=1u
M10368 net3113 n4251 VDD VDD pmos w=2u l=1u
M10369 n4296 n4249 VDD VDD pmos w=2u l=1u
M10370 n4296 n4249 VSS VSS nmos w=1u l=1u
M10371 n4243 n4299 VSS VSS nmos w=1u l=1u
M10372 n4243 n4298 VSS VSS nmos w=1u l=1u
M10373 n4243 n4299 net3114 VDD pmos w=2u l=1u
M10374 net3114 n4298 VDD VDD pmos w=2u l=1u
M10375 n4299 net3115 VSS VSS nmos w=1u l=1u
M10376 net3116 n4240 VSS VSS nmos w=1u l=1u
M10377 net3115 n4241 net3116 VSS nmos w=1u l=1u
M10378 net3115 n4240 VDD VDD pmos w=2u l=1u
M10379 net3115 n4241 VDD VDD pmos w=2u l=1u
M10380 n4299 net3115 VDD VDD pmos w=2u l=1u
M10381 n4298 n4239 VDD VDD pmos w=2u l=1u
M10382 n4298 n4239 VSS VSS nmos w=1u l=1u
M10383 n4233 n4301 VSS VSS nmos w=1u l=1u
M10384 n4233 n4300 VSS VSS nmos w=1u l=1u
M10385 n4233 n4301 net3117 VDD pmos w=2u l=1u
M10386 net3117 n4300 VDD VDD pmos w=2u l=1u
M10387 n4301 net3118 VSS VSS nmos w=1u l=1u
M10388 net3119 n4230 VSS VSS nmos w=1u l=1u
M10389 net3118 n4231 net3119 VSS nmos w=1u l=1u
M10390 net3118 n4230 VDD VDD pmos w=2u l=1u
M10391 net3118 n4231 VDD VDD pmos w=2u l=1u
M10392 n4301 net3118 VDD VDD pmos w=2u l=1u
M10393 n4300 n4229 VDD VDD pmos w=2u l=1u
M10394 n4300 n4229 VSS VSS nmos w=1u l=1u
M10395 n4223 n4303 VSS VSS nmos w=1u l=1u
M10396 n4223 n4302 VSS VSS nmos w=1u l=1u
M10397 n4223 n4303 net3120 VDD pmos w=2u l=1u
M10398 net3120 n4302 VDD VDD pmos w=2u l=1u
M10399 n4303 n4305 VSS VSS nmos w=1u l=1u
M10400 n4303 n4304 VSS VSS nmos w=1u l=1u
M10401 n4303 n4305 net3121 VDD pmos w=2u l=1u
M10402 net3121 n4304 VDD VDD pmos w=2u l=1u
M10403 n4304 n4221 VDD VDD pmos w=2u l=1u
M10404 n4304 n4221 VSS VSS nmos w=1u l=1u
M10405 n4302 n4219 VDD VDD pmos w=2u l=1u
M10406 n4302 n4219 VSS VSS nmos w=1u l=1u
M10407 n4213 n4307 VSS VSS nmos w=1u l=1u
M10408 n4213 n4306 VSS VSS nmos w=1u l=1u
M10409 n4213 n4307 net3122 VDD pmos w=2u l=1u
M10410 net3122 n4306 VDD VDD pmos w=2u l=1u
M10411 n4307 n4309 VSS VSS nmos w=1u l=1u
M10412 n4307 n4308 VSS VSS nmos w=1u l=1u
M10413 n4307 n4309 net3123 VDD pmos w=2u l=1u
M10414 net3123 n4308 VDD VDD pmos w=2u l=1u
M10415 n4308 n4212 VDD VDD pmos w=2u l=1u
M10416 n4308 n4212 VSS VSS nmos w=1u l=1u
M10417 n4306 n4210 VDD VDD pmos w=2u l=1u
M10418 n4306 n4210 VSS VSS nmos w=1u l=1u
M10419 n4204 n4311 VSS VSS nmos w=1u l=1u
M10420 n4204 n4310 VSS VSS nmos w=1u l=1u
M10421 n4204 n4311 net3124 VDD pmos w=2u l=1u
M10422 net3124 n4310 VDD VDD pmos w=2u l=1u
M10423 n4311 n4202 VSS VSS nmos w=1u l=1u
M10424 n4311 n4203 VSS VSS nmos w=1u l=1u
M10425 n4311 n4202 net3125 VDD pmos w=2u l=1u
M10426 net3125 n4203 VDD VDD pmos w=2u l=1u
M10427 n4310 n4201 VDD VDD pmos w=2u l=1u
M10428 n4310 n4201 VSS VSS nmos w=1u l=1u
M10429 net3126 n4203 VSS VSS nmos w=1u l=1u
M10430 net3127 n4312 VSS VSS nmos w=1u l=1u
M10431 N4591 net3128 VSS VSS nmos w=1u l=1u
M10432 net3128 n4203 net3129 VSS nmos w=1u l=1u
M10433 net3128 net3126 net3127 VSS nmos w=1u l=1u
M10434 net3129 net3127 VSS VSS nmos w=1u l=1u
M10435 net3128 net3126 net3130 VDD pmos w=2u l=1u
M10436 net3126 n4203 VDD VDD pmos w=2u l=1u
M10437 net3127 n4203 net3128 VDD pmos w=2u l=1u
M10438 net3127 n4312 VDD VDD pmos w=2u l=1u
M10439 N4591 net3128 VDD VDD pmos w=2u l=1u
M10440 net3130 net3127 VDD VDD pmos w=2u l=1u
M10441 n4203 n2445 VSS VSS nmos w=1u l=1u
M10442 n4203 n3929 VSS VSS nmos w=1u l=1u
M10443 n4203 n2445 net3131 VDD pmos w=2u l=1u
M10444 net3131 n3929 VDD VDD pmos w=2u l=1u
M10445 n2445 N443 VDD VDD pmos w=2u l=1u
M10446 n2445 N443 VSS VSS nmos w=1u l=1u
M10447 n4312 n4202 VDD VDD pmos w=2u l=1u
M10448 n4312 n4202 VSS VSS nmos w=1u l=1u
M10449 n4202 n4201 net3132 VSS nmos w=1u l=1u
M10450 net3132 n4313 VSS VSS nmos w=1u l=1u
M10451 n4202 n4201 VDD VDD pmos w=2u l=1u
M10452 n4202 n4313 VDD VDD pmos w=2u l=1u
M10453 n4201 n4315 net3133 VSS nmos w=1u l=1u
M10454 net3133 n4314 VSS VSS nmos w=1u l=1u
M10455 n4201 n4315 VDD VDD pmos w=2u l=1u
M10456 n4201 n4314 VDD VDD pmos w=2u l=1u
M10457 n4315 n4317 net3134 VSS nmos w=1u l=1u
M10458 net3134 n4316 VSS VSS nmos w=1u l=1u
M10459 n4315 n4317 VDD VDD pmos w=2u l=1u
M10460 n4315 n4316 VDD VDD pmos w=2u l=1u
M10461 n4316 net3135 VSS VSS nmos w=1u l=1u
M10462 net3135 n4318 VSS VSS nmos w=1u l=1u
M10463 net3135 n4319 VSS VSS nmos w=1u l=1u
M10464 net3135 n4319 net3136 VDD pmos w=2u l=1u
M10465 n4316 net3135 VDD VDD pmos w=2u l=1u
M10466 net3136 n4318 VDD VDD pmos w=2u l=1u
M10467 net3137 n4211 VSS VSS nmos w=1u l=1u
M10468 net3138 n4212 VSS VSS nmos w=1u l=1u
M10469 n4314 net3139 VSS VSS nmos w=1u l=1u
M10470 net3139 n4211 net3140 VSS nmos w=1u l=1u
M10471 net3139 net3137 net3138 VSS nmos w=1u l=1u
M10472 net3140 net3138 VSS VSS nmos w=1u l=1u
M10473 net3139 net3137 net3141 VDD pmos w=2u l=1u
M10474 net3137 n4211 VDD VDD pmos w=2u l=1u
M10475 net3138 n4211 net3139 VDD pmos w=2u l=1u
M10476 net3138 n4212 VDD VDD pmos w=2u l=1u
M10477 n4314 net3139 VDD VDD pmos w=2u l=1u
M10478 net3141 net3138 VDD VDD pmos w=2u l=1u
M10479 n4211 n4309 VDD VDD pmos w=2u l=1u
M10480 n4211 n4309 VSS VSS nmos w=1u l=1u
M10481 n4313 n4321 net3142 VSS nmos w=1u l=1u
M10482 net3142 n4320 VSS VSS nmos w=1u l=1u
M10483 n4313 n4321 VDD VDD pmos w=2u l=1u
M10484 n4313 n4320 VDD VDD pmos w=2u l=1u
M10485 net3143 n4212 VSS VSS nmos w=1u l=1u
M10486 net3144 n4309 VSS VSS nmos w=1u l=1u
M10487 n4321 net3145 VSS VSS nmos w=1u l=1u
M10488 net3145 n4212 net3146 VSS nmos w=1u l=1u
M10489 net3145 net3143 net3144 VSS nmos w=1u l=1u
M10490 net3146 net3144 VSS VSS nmos w=1u l=1u
M10491 net3145 net3143 net3147 VDD pmos w=2u l=1u
M10492 net3143 n4212 VDD VDD pmos w=2u l=1u
M10493 net3144 n4212 net3145 VDD pmos w=2u l=1u
M10494 net3144 n4309 VDD VDD pmos w=2u l=1u
M10495 n4321 net3145 VDD VDD pmos w=2u l=1u
M10496 net3147 net3144 VDD VDD pmos w=2u l=1u
M10497 n4212 N426 net3148 VSS nmos w=1u l=1u
M10498 net3148 N18 VSS VSS nmos w=1u l=1u
M10499 n4212 N426 VDD VDD pmos w=2u l=1u
M10500 n4212 N18 VDD VDD pmos w=2u l=1u
M10501 n4309 n4210 net3149 VSS nmos w=1u l=1u
M10502 net3149 n4322 VSS VSS nmos w=1u l=1u
M10503 n4309 n4210 VDD VDD pmos w=2u l=1u
M10504 n4309 n4322 VDD VDD pmos w=2u l=1u
M10505 n4210 n4324 net3150 VSS nmos w=1u l=1u
M10506 net3150 n4323 VSS VSS nmos w=1u l=1u
M10507 n4210 n4324 VDD VDD pmos w=2u l=1u
M10508 n4210 n4323 VDD VDD pmos w=2u l=1u
M10509 n4324 n4326 net3151 VSS nmos w=1u l=1u
M10510 net3151 n4325 VSS VSS nmos w=1u l=1u
M10511 n4324 n4326 VDD VDD pmos w=2u l=1u
M10512 n4324 n4325 VDD VDD pmos w=2u l=1u
M10513 n4325 n4328 net3152 VSS nmos w=1u l=1u
M10514 net3152 n4327 VSS VSS nmos w=1u l=1u
M10515 n4325 n4328 VDD VDD pmos w=2u l=1u
M10516 n4325 n4327 VDD VDD pmos w=2u l=1u
M10517 net3153 n4220 VSS VSS nmos w=1u l=1u
M10518 net3154 n4221 VSS VSS nmos w=1u l=1u
M10519 n4323 net3155 VSS VSS nmos w=1u l=1u
M10520 net3155 n4220 net3156 VSS nmos w=1u l=1u
M10521 net3155 net3153 net3154 VSS nmos w=1u l=1u
M10522 net3156 net3154 VSS VSS nmos w=1u l=1u
M10523 net3155 net3153 net3157 VDD pmos w=2u l=1u
M10524 net3153 n4220 VDD VDD pmos w=2u l=1u
M10525 net3154 n4220 net3155 VDD pmos w=2u l=1u
M10526 net3154 n4221 VDD VDD pmos w=2u l=1u
M10527 n4323 net3155 VDD VDD pmos w=2u l=1u
M10528 net3157 net3154 VDD VDD pmos w=2u l=1u
M10529 n4220 n4305 VDD VDD pmos w=2u l=1u
M10530 n4220 n4305 VSS VSS nmos w=1u l=1u
M10531 n4322 n4330 net3158 VSS nmos w=1u l=1u
M10532 net3158 n4329 VSS VSS nmos w=1u l=1u
M10533 n4322 n4330 VDD VDD pmos w=2u l=1u
M10534 n4322 n4329 VDD VDD pmos w=2u l=1u
M10535 net3159 n4221 VSS VSS nmos w=1u l=1u
M10536 net3160 n4305 VSS VSS nmos w=1u l=1u
M10537 n4330 net3161 VSS VSS nmos w=1u l=1u
M10538 net3161 n4221 net3162 VSS nmos w=1u l=1u
M10539 net3161 net3159 net3160 VSS nmos w=1u l=1u
M10540 net3162 net3160 VSS VSS nmos w=1u l=1u
M10541 net3161 net3159 net3163 VDD pmos w=2u l=1u
M10542 net3159 n4221 VDD VDD pmos w=2u l=1u
M10543 net3160 n4221 net3161 VDD pmos w=2u l=1u
M10544 net3160 n4305 VDD VDD pmos w=2u l=1u
M10545 n4330 net3161 VDD VDD pmos w=2u l=1u
M10546 net3163 net3160 VDD VDD pmos w=2u l=1u
M10547 n4221 N409 net3164 VSS nmos w=1u l=1u
M10548 net3164 N35 VSS VSS nmos w=1u l=1u
M10549 n4221 N409 VDD VDD pmos w=2u l=1u
M10550 n4221 N35 VDD VDD pmos w=2u l=1u
M10551 n4305 n4219 net3165 VSS nmos w=1u l=1u
M10552 net3165 n4331 VSS VSS nmos w=1u l=1u
M10553 n4305 n4219 VDD VDD pmos w=2u l=1u
M10554 n4305 n4331 VDD VDD pmos w=2u l=1u
M10555 n4219 n4333 net3166 VSS nmos w=1u l=1u
M10556 net3166 n4332 VSS VSS nmos w=1u l=1u
M10557 n4219 n4333 VDD VDD pmos w=2u l=1u
M10558 n4219 n4332 VDD VDD pmos w=2u l=1u
M10559 n4333 n4335 net3167 VSS nmos w=1u l=1u
M10560 net3167 n4334 VSS VSS nmos w=1u l=1u
M10561 n4333 n4335 VDD VDD pmos w=2u l=1u
M10562 n4333 n4334 VDD VDD pmos w=2u l=1u
M10563 n4334 n4337 net3168 VSS nmos w=1u l=1u
M10564 net3168 n4336 VSS VSS nmos w=1u l=1u
M10565 n4334 n4337 VDD VDD pmos w=2u l=1u
M10566 n4334 n4336 VDD VDD pmos w=2u l=1u
M10567 net3169 n4230 VSS VSS nmos w=1u l=1u
M10568 net3170 n4231 VSS VSS nmos w=1u l=1u
M10569 n4332 net3171 VSS VSS nmos w=1u l=1u
M10570 net3171 n4230 net3172 VSS nmos w=1u l=1u
M10571 net3171 net3169 net3170 VSS nmos w=1u l=1u
M10572 net3172 net3170 VSS VSS nmos w=1u l=1u
M10573 net3171 net3169 net3173 VDD pmos w=2u l=1u
M10574 net3169 n4230 VDD VDD pmos w=2u l=1u
M10575 net3170 n4230 net3171 VDD pmos w=2u l=1u
M10576 net3170 n4231 VDD VDD pmos w=2u l=1u
M10577 n4332 net3171 VDD VDD pmos w=2u l=1u
M10578 net3173 net3170 VDD VDD pmos w=2u l=1u
M10579 n4230 n4338 VDD VDD pmos w=2u l=1u
M10580 n4230 n4338 VSS VSS nmos w=1u l=1u
M10581 n4331 n4340 net3174 VSS nmos w=1u l=1u
M10582 net3174 n4339 VSS VSS nmos w=1u l=1u
M10583 n4331 n4340 VDD VDD pmos w=2u l=1u
M10584 n4331 n4339 VDD VDD pmos w=2u l=1u
M10585 net3175 n4231 VSS VSS nmos w=1u l=1u
M10586 net3176 n4338 VSS VSS nmos w=1u l=1u
M10587 n4340 net3177 VSS VSS nmos w=1u l=1u
M10588 net3177 n4231 net3178 VSS nmos w=1u l=1u
M10589 net3177 net3175 net3176 VSS nmos w=1u l=1u
M10590 net3178 net3176 VSS VSS nmos w=1u l=1u
M10591 net3177 net3175 net3179 VDD pmos w=2u l=1u
M10592 net3175 n4231 VDD VDD pmos w=2u l=1u
M10593 net3176 n4231 net3177 VDD pmos w=2u l=1u
M10594 net3176 n4338 VDD VDD pmos w=2u l=1u
M10595 n4340 net3177 VDD VDD pmos w=2u l=1u
M10596 net3179 net3176 VDD VDD pmos w=2u l=1u
M10597 n4231 N392 net3180 VSS nmos w=1u l=1u
M10598 net3180 N52 VSS VSS nmos w=1u l=1u
M10599 n4231 N392 VDD VDD pmos w=2u l=1u
M10600 n4231 N52 VDD VDD pmos w=2u l=1u
M10601 n4338 n4229 net3181 VSS nmos w=1u l=1u
M10602 net3181 n4341 VSS VSS nmos w=1u l=1u
M10603 n4338 n4229 VDD VDD pmos w=2u l=1u
M10604 n4338 n4341 VDD VDD pmos w=2u l=1u
M10605 n4229 n4343 net3182 VSS nmos w=1u l=1u
M10606 net3182 n4342 VSS VSS nmos w=1u l=1u
M10607 n4229 n4343 VDD VDD pmos w=2u l=1u
M10608 n4229 n4342 VDD VDD pmos w=2u l=1u
M10609 n4343 n4345 net3183 VSS nmos w=1u l=1u
M10610 net3183 n4344 VSS VSS nmos w=1u l=1u
M10611 n4343 n4345 VDD VDD pmos w=2u l=1u
M10612 n4343 n4344 VDD VDD pmos w=2u l=1u
M10613 n4344 n4347 net3184 VSS nmos w=1u l=1u
M10614 net3184 n4346 VSS VSS nmos w=1u l=1u
M10615 n4344 n4347 VDD VDD pmos w=2u l=1u
M10616 n4344 n4346 VDD VDD pmos w=2u l=1u
M10617 net3185 n4240 VSS VSS nmos w=1u l=1u
M10618 net3186 n4241 VSS VSS nmos w=1u l=1u
M10619 n4342 net3187 VSS VSS nmos w=1u l=1u
M10620 net3187 n4240 net3188 VSS nmos w=1u l=1u
M10621 net3187 net3185 net3186 VSS nmos w=1u l=1u
M10622 net3188 net3186 VSS VSS nmos w=1u l=1u
M10623 net3187 net3185 net3189 VDD pmos w=2u l=1u
M10624 net3185 n4240 VDD VDD pmos w=2u l=1u
M10625 net3186 n4240 net3187 VDD pmos w=2u l=1u
M10626 net3186 n4241 VDD VDD pmos w=2u l=1u
M10627 n4342 net3187 VDD VDD pmos w=2u l=1u
M10628 net3189 net3186 VDD VDD pmos w=2u l=1u
M10629 n4240 n4348 VDD VDD pmos w=2u l=1u
M10630 n4240 n4348 VSS VSS nmos w=1u l=1u
M10631 n4341 n4350 net3190 VSS nmos w=1u l=1u
M10632 net3190 n4349 VSS VSS nmos w=1u l=1u
M10633 n4341 n4350 VDD VDD pmos w=2u l=1u
M10634 n4341 n4349 VDD VDD pmos w=2u l=1u
M10635 net3191 n4241 VSS VSS nmos w=1u l=1u
M10636 net3192 n4348 VSS VSS nmos w=1u l=1u
M10637 n4350 net3193 VSS VSS nmos w=1u l=1u
M10638 net3193 n4241 net3194 VSS nmos w=1u l=1u
M10639 net3193 net3191 net3192 VSS nmos w=1u l=1u
M10640 net3194 net3192 VSS VSS nmos w=1u l=1u
M10641 net3193 net3191 net3195 VDD pmos w=2u l=1u
M10642 net3191 n4241 VDD VDD pmos w=2u l=1u
M10643 net3192 n4241 net3193 VDD pmos w=2u l=1u
M10644 net3192 n4348 VDD VDD pmos w=2u l=1u
M10645 n4350 net3193 VDD VDD pmos w=2u l=1u
M10646 net3195 net3192 VDD VDD pmos w=2u l=1u
M10647 n4241 N375 net3196 VSS nmos w=1u l=1u
M10648 net3196 N69 VSS VSS nmos w=1u l=1u
M10649 n4241 N375 VDD VDD pmos w=2u l=1u
M10650 n4241 N69 VDD VDD pmos w=2u l=1u
M10651 n4348 n4239 net3197 VSS nmos w=1u l=1u
M10652 net3197 n4351 VSS VSS nmos w=1u l=1u
M10653 n4348 n4239 VDD VDD pmos w=2u l=1u
M10654 n4348 n4351 VDD VDD pmos w=2u l=1u
M10655 n4239 n4353 net3198 VSS nmos w=1u l=1u
M10656 net3198 n4352 VSS VSS nmos w=1u l=1u
M10657 n4239 n4353 VDD VDD pmos w=2u l=1u
M10658 n4239 n4352 VDD VDD pmos w=2u l=1u
M10659 n4353 n4355 net3199 VSS nmos w=1u l=1u
M10660 net3199 n4354 VSS VSS nmos w=1u l=1u
M10661 n4353 n4355 VDD VDD pmos w=2u l=1u
M10662 n4353 n4354 VDD VDD pmos w=2u l=1u
M10663 n4354 net3200 VSS VSS nmos w=1u l=1u
M10664 net3200 n4356 VSS VSS nmos w=1u l=1u
M10665 net3200 n4357 VSS VSS nmos w=1u l=1u
M10666 net3200 n4357 net3201 VDD pmos w=2u l=1u
M10667 n4354 net3200 VDD VDD pmos w=2u l=1u
M10668 net3201 n4356 VDD VDD pmos w=2u l=1u
M10669 net3202 n4250 VSS VSS nmos w=1u l=1u
M10670 net3203 n4251 VSS VSS nmos w=1u l=1u
M10671 n4352 net3204 VSS VSS nmos w=1u l=1u
M10672 net3204 n4250 net3205 VSS nmos w=1u l=1u
M10673 net3204 net3202 net3203 VSS nmos w=1u l=1u
M10674 net3205 net3203 VSS VSS nmos w=1u l=1u
M10675 net3204 net3202 net3206 VDD pmos w=2u l=1u
M10676 net3202 n4250 VDD VDD pmos w=2u l=1u
M10677 net3203 n4250 net3204 VDD pmos w=2u l=1u
M10678 net3203 n4251 VDD VDD pmos w=2u l=1u
M10679 n4352 net3204 VDD VDD pmos w=2u l=1u
M10680 net3206 net3203 VDD VDD pmos w=2u l=1u
M10681 n4251 n4358 VDD VDD pmos w=2u l=1u
M10682 n4251 n4358 VSS VSS nmos w=1u l=1u
M10683 n4351 n4360 net3207 VSS nmos w=1u l=1u
M10684 net3207 n4359 VSS VSS nmos w=1u l=1u
M10685 n4351 n4360 VDD VDD pmos w=2u l=1u
M10686 n4351 n4359 VDD VDD pmos w=2u l=1u
M10687 net3208 n4358 VSS VSS nmos w=1u l=1u
M10688 net3209 n4250 VSS VSS nmos w=1u l=1u
M10689 n4360 net3210 VSS VSS nmos w=1u l=1u
M10690 net3210 n4358 net3211 VSS nmos w=1u l=1u
M10691 net3210 net3208 net3209 VSS nmos w=1u l=1u
M10692 net3211 net3209 VSS VSS nmos w=1u l=1u
M10693 net3210 net3208 net3212 VDD pmos w=2u l=1u
M10694 net3208 n4358 VDD VDD pmos w=2u l=1u
M10695 net3209 n4358 net3210 VDD pmos w=2u l=1u
M10696 net3209 n4250 VDD VDD pmos w=2u l=1u
M10697 n4360 net3210 VDD VDD pmos w=2u l=1u
M10698 net3212 net3209 VDD VDD pmos w=2u l=1u
M10699 n4358 N358 net3213 VSS nmos w=1u l=1u
M10700 net3213 N86 VSS VSS nmos w=1u l=1u
M10701 n4358 N358 VDD VDD pmos w=2u l=1u
M10702 n4358 N86 VDD VDD pmos w=2u l=1u
M10703 n4250 n4249 net3214 VSS nmos w=1u l=1u
M10704 net3214 n4361 VSS VSS nmos w=1u l=1u
M10705 n4250 n4249 VDD VDD pmos w=2u l=1u
M10706 n4250 n4361 VDD VDD pmos w=2u l=1u
M10707 n4249 n4363 net3215 VSS nmos w=1u l=1u
M10708 net3215 n4362 VSS VSS nmos w=1u l=1u
M10709 n4249 n4363 VDD VDD pmos w=2u l=1u
M10710 n4249 n4362 VDD VDD pmos w=2u l=1u
M10711 n4363 n4365 net3216 VSS nmos w=1u l=1u
M10712 net3216 n4364 VSS VSS nmos w=1u l=1u
M10713 n4363 n4365 VDD VDD pmos w=2u l=1u
M10714 n4363 n4364 VDD VDD pmos w=2u l=1u
M10715 n4364 n4367 net3217 VSS nmos w=1u l=1u
M10716 net3217 n4366 VSS VSS nmos w=1u l=1u
M10717 n4364 n4367 VDD VDD pmos w=2u l=1u
M10718 n4364 n4366 VDD VDD pmos w=2u l=1u
M10719 net3218 n4260 VSS VSS nmos w=1u l=1u
M10720 net3219 n4261 VSS VSS nmos w=1u l=1u
M10721 n4362 net3220 VSS VSS nmos w=1u l=1u
M10722 net3220 n4260 net3221 VSS nmos w=1u l=1u
M10723 net3220 net3218 net3219 VSS nmos w=1u l=1u
M10724 net3221 net3219 VSS VSS nmos w=1u l=1u
M10725 net3220 net3218 net3222 VDD pmos w=2u l=1u
M10726 net3218 n4260 VDD VDD pmos w=2u l=1u
M10727 net3219 n4260 net3220 VDD pmos w=2u l=1u
M10728 net3219 n4261 VDD VDD pmos w=2u l=1u
M10729 n4362 net3220 VDD VDD pmos w=2u l=1u
M10730 net3222 net3219 VDD VDD pmos w=2u l=1u
M10731 n4260 n4368 VDD VDD pmos w=2u l=1u
M10732 n4260 n4368 VSS VSS nmos w=1u l=1u
M10733 n4361 n4370 net3223 VSS nmos w=1u l=1u
M10734 net3223 n4369 VSS VSS nmos w=1u l=1u
M10735 n4361 n4370 VDD VDD pmos w=2u l=1u
M10736 n4361 n4369 VDD VDD pmos w=2u l=1u
M10737 net3224 n4261 VSS VSS nmos w=1u l=1u
M10738 net3225 n4368 VSS VSS nmos w=1u l=1u
M10739 n4370 net3226 VSS VSS nmos w=1u l=1u
M10740 net3226 n4261 net3227 VSS nmos w=1u l=1u
M10741 net3226 net3224 net3225 VSS nmos w=1u l=1u
M10742 net3227 net3225 VSS VSS nmos w=1u l=1u
M10743 net3226 net3224 net3228 VDD pmos w=2u l=1u
M10744 net3224 n4261 VDD VDD pmos w=2u l=1u
M10745 net3225 n4261 net3226 VDD pmos w=2u l=1u
M10746 net3225 n4368 VDD VDD pmos w=2u l=1u
M10747 n4370 net3226 VDD VDD pmos w=2u l=1u
M10748 net3228 net3225 VDD VDD pmos w=2u l=1u
M10749 n4261 N341 net3229 VSS nmos w=1u l=1u
M10750 net3229 N103 VSS VSS nmos w=1u l=1u
M10751 n4261 N341 VDD VDD pmos w=2u l=1u
M10752 n4261 N103 VDD VDD pmos w=2u l=1u
M10753 n4368 n4259 net3230 VSS nmos w=1u l=1u
M10754 net3230 n4371 VSS VSS nmos w=1u l=1u
M10755 n4368 n4259 VDD VDD pmos w=2u l=1u
M10756 n4368 n4371 VDD VDD pmos w=2u l=1u
M10757 n4259 n4373 net3231 VSS nmos w=1u l=1u
M10758 net3231 n4372 VSS VSS nmos w=1u l=1u
M10759 n4259 n4373 VDD VDD pmos w=2u l=1u
M10760 n4259 n4372 VDD VDD pmos w=2u l=1u
M10761 n4373 net3232 VSS VSS nmos w=1u l=1u
M10762 net3232 n4374 VSS VSS nmos w=1u l=1u
M10763 net3232 n4375 VSS VSS nmos w=1u l=1u
M10764 net3232 n4375 net3233 VDD pmos w=2u l=1u
M10765 n4373 net3232 VDD VDD pmos w=2u l=1u
M10766 net3233 n4374 VDD VDD pmos w=2u l=1u
M10767 n4372 net3234 VSS VSS nmos w=1u l=1u
M10768 net3235 n4376 VSS VSS nmos w=1u l=1u
M10769 net3234 n4293 net3235 VSS nmos w=1u l=1u
M10770 net3234 n4376 VDD VDD pmos w=2u l=1u
M10771 net3234 n4293 VDD VDD pmos w=2u l=1u
M10772 n4372 net3234 VDD VDD pmos w=2u l=1u
M10773 n4371 n4378 net3236 VSS nmos w=1u l=1u
M10774 net3236 n4377 VSS VSS nmos w=1u l=1u
M10775 n4371 n4378 VDD VDD pmos w=2u l=1u
M10776 n4371 n4377 VDD VDD pmos w=2u l=1u
M10777 n4378 n4293 net3237 VSS nmos w=1u l=1u
M10778 net3237 n4376 VSS VSS nmos w=1u l=1u
M10779 n4378 n4293 VDD VDD pmos w=2u l=1u
M10780 n4378 n4376 VDD VDD pmos w=2u l=1u
M10781 n4293 n4380 net3238 VSS nmos w=1u l=1u
M10782 net3238 n4379 VSS VSS nmos w=1u l=1u
M10783 n4293 n4380 VDD VDD pmos w=2u l=1u
M10784 n4293 n4379 VDD VDD pmos w=2u l=1u
M10785 n4380 N324 net3239 VSS nmos w=1u l=1u
M10786 net3239 N120 VSS VSS nmos w=1u l=1u
M10787 n4380 N324 VDD VDD pmos w=2u l=1u
M10788 n4380 N120 VDD VDD pmos w=2u l=1u
M10789 n4376 N120 net3240 VSS nmos w=1u l=1u
M10790 net3240 n4381 VSS VSS nmos w=1u l=1u
M10791 n4376 N120 VDD VDD pmos w=2u l=1u
M10792 n4376 n4381 VDD VDD pmos w=2u l=1u
M10793 n4381 n3257 VSS VSS nmos w=1u l=1u
M10794 n4381 n4379 VSS VSS nmos w=1u l=1u
M10795 n4381 n3257 net3241 VDD pmos w=2u l=1u
M10796 net3241 n4379 VDD VDD pmos w=2u l=1u
M10797 n4379 n4269 VSS VSS nmos w=1u l=1u
M10798 n4379 n4382 VSS VSS nmos w=1u l=1u
M10799 n4379 n4269 net3242 VDD pmos w=2u l=1u
M10800 net3242 n4382 VDD VDD pmos w=2u l=1u
M10801 n4269 n4384 VSS VSS nmos w=1u l=1u
M10802 n4269 n4383 VSS VSS nmos w=1u l=1u
M10803 n4269 n4384 net3243 VDD pmos w=2u l=1u
M10804 net3243 n4383 VDD VDD pmos w=2u l=1u
M10805 n4382 net3244 VSS VSS nmos w=1u l=1u
M10806 net3245 n4383 VSS VSS nmos w=1u l=1u
M10807 net3244 n4384 net3245 VSS nmos w=1u l=1u
M10808 net3244 n4383 VDD VDD pmos w=2u l=1u
M10809 net3244 n4384 VDD VDD pmos w=2u l=1u
M10810 n4382 net3244 VDD VDD pmos w=2u l=1u
M10811 n4383 n4385 net3246 VSS nmos w=1u l=1u
M10812 net3246 n4291 VSS VSS nmos w=1u l=1u
M10813 n4383 n4385 VDD VDD pmos w=2u l=1u
M10814 n4383 n4291 VDD VDD pmos w=2u l=1u
M10815 n4385 N137 net3247 VSS nmos w=1u l=1u
M10816 net3247 n4386 VSS VSS nmos w=1u l=1u
M10817 n4385 N137 VDD VDD pmos w=2u l=1u
M10818 n4385 n4386 VDD VDD pmos w=2u l=1u
M10819 n4386 n3411 VSS VSS nmos w=1u l=1u
M10820 n4386 n4387 VSS VSS nmos w=1u l=1u
M10821 n4386 n3411 net3248 VDD pmos w=2u l=1u
M10822 net3248 n4387 VDD VDD pmos w=2u l=1u
M10823 n4291 n4388 net3249 VSS nmos w=1u l=1u
M10824 net3249 n4387 VSS VSS nmos w=1u l=1u
M10825 n4291 n4388 VDD VDD pmos w=2u l=1u
M10826 n4291 n4387 VDD VDD pmos w=2u l=1u
M10827 n4388 N307 net3250 VSS nmos w=1u l=1u
M10828 net3250 N137 VSS VSS nmos w=1u l=1u
M10829 n4388 N307 VDD VDD pmos w=2u l=1u
M10830 n4388 N137 VDD VDD pmos w=2u l=1u
M10831 n4387 net3251 VSS VSS nmos w=1u l=1u
M10832 net3252 n4389 VSS VSS nmos w=1u l=1u
M10833 net3251 n4292 net3252 VSS nmos w=1u l=1u
M10834 net3251 n4389 VDD VDD pmos w=2u l=1u
M10835 net3251 n4292 VDD VDD pmos w=2u l=1u
M10836 n4387 net3251 VDD VDD pmos w=2u l=1u
M10837 n4389 net3253 VSS VSS nmos w=1u l=1u
M10838 net3253 n4390 VSS VSS nmos w=1u l=1u
M10839 net3253 n4284 VSS VSS nmos w=1u l=1u
M10840 net3253 n4284 net3254 VDD pmos w=2u l=1u
M10841 n4389 net3253 VDD VDD pmos w=2u l=1u
M10842 net3254 n4390 VDD VDD pmos w=2u l=1u
M10843 n4284 n4285 VDD VDD pmos w=2u l=1u
M10844 n4284 n4285 VSS VSS nmos w=1u l=1u
M10845 n4292 n4391 net3255 VSS nmos w=1u l=1u
M10846 net3255 n4390 VSS VSS nmos w=1u l=1u
M10847 n4292 n4391 VDD VDD pmos w=2u l=1u
M10848 n4292 n4390 VDD VDD pmos w=2u l=1u
M10849 n4391 n4285 net3256 VSS nmos w=1u l=1u
M10850 net3256 n4392 VSS VSS nmos w=1u l=1u
M10851 n4391 n4285 VDD VDD pmos w=2u l=1u
M10852 n4391 n4392 VDD VDD pmos w=2u l=1u
M10853 n4285 N171 net3257 VSS nmos w=1u l=1u
M10854 net3257 n4393 VSS VSS nmos w=1u l=1u
M10855 n4285 N171 VDD VDD pmos w=2u l=1u
M10856 n4285 n4393 VDD VDD pmos w=2u l=1u
M10857 n4393 net3258 VSS VSS nmos w=1u l=1u
M10858 net3259 N154 VSS VSS nmos w=1u l=1u
M10859 net3258 n3741 net3259 VSS nmos w=1u l=1u
M10860 net3258 N154 VDD VDD pmos w=2u l=1u
M10861 net3258 n3741 VDD VDD pmos w=2u l=1u
M10862 n4393 net3258 VDD VDD pmos w=2u l=1u
M10863 n4392 n4395 net3260 VSS nmos w=1u l=1u
M10864 net3260 n4394 VSS VSS nmos w=1u l=1u
M10865 n4392 n4395 VDD VDD pmos w=2u l=1u
M10866 n4392 n4394 VDD VDD pmos w=2u l=1u
M10867 n4395 N273 net3261 VSS nmos w=1u l=1u
M10868 net3261 N171 VSS VSS nmos w=1u l=1u
M10869 n4395 N273 VDD VDD pmos w=2u l=1u
M10870 n4395 N171 VDD VDD pmos w=2u l=1u
M10871 n4394 N290 net3262 VSS nmos w=1u l=1u
M10872 net3262 N154 VSS VSS nmos w=1u l=1u
M10873 n4394 N290 VDD VDD pmos w=2u l=1u
M10874 n4394 N154 VDD VDD pmos w=2u l=1u
M10875 n4384 net3263 VSS VSS nmos w=1u l=1u
M10876 net3264 n4397 VSS VSS nmos w=1u l=1u
M10877 net3263 n4396 net3264 VSS nmos w=1u l=1u
M10878 net3263 n4397 VDD VDD pmos w=2u l=1u
M10879 net3263 n4396 VDD VDD pmos w=2u l=1u
M10880 n4384 net3263 VDD VDD pmos w=2u l=1u
M10881 n4377 n4374 VSS VSS nmos w=1u l=1u
M10882 n4377 n4375 VSS VSS nmos w=1u l=1u
M10883 n4377 n4374 net3265 VDD pmos w=2u l=1u
M10884 net3265 n4375 VDD VDD pmos w=2u l=1u
M10885 n4374 n4398 VDD VDD pmos w=2u l=1u
M10886 n4374 n4398 VSS VSS nmos w=1u l=1u
M10887 n4369 n4400 VSS VSS nmos w=1u l=1u
M10888 n4369 n4399 VSS VSS nmos w=1u l=1u
M10889 n4369 n4400 net3266 VDD pmos w=2u l=1u
M10890 net3266 n4399 VDD VDD pmos w=2u l=1u
M10891 n4400 net3267 VSS VSS nmos w=1u l=1u
M10892 net3268 n4366 VSS VSS nmos w=1u l=1u
M10893 net3267 n4367 net3268 VSS nmos w=1u l=1u
M10894 net3267 n4366 VDD VDD pmos w=2u l=1u
M10895 net3267 n4367 VDD VDD pmos w=2u l=1u
M10896 n4400 net3267 VDD VDD pmos w=2u l=1u
M10897 n4399 n4365 VDD VDD pmos w=2u l=1u
M10898 n4399 n4365 VSS VSS nmos w=1u l=1u
M10899 n4359 n4402 VSS VSS nmos w=1u l=1u
M10900 n4359 n4401 VSS VSS nmos w=1u l=1u
M10901 n4359 n4402 net3269 VDD pmos w=2u l=1u
M10902 net3269 n4401 VDD VDD pmos w=2u l=1u
M10903 n4402 n4356 VSS VSS nmos w=1u l=1u
M10904 n4402 n4357 VSS VSS nmos w=1u l=1u
M10905 n4402 n4356 net3270 VDD pmos w=2u l=1u
M10906 net3270 n4357 VDD VDD pmos w=2u l=1u
M10907 n4401 n4355 VDD VDD pmos w=2u l=1u
M10908 n4401 n4355 VSS VSS nmos w=1u l=1u
M10909 n4349 n4404 VSS VSS nmos w=1u l=1u
M10910 n4349 n4403 VSS VSS nmos w=1u l=1u
M10911 n4349 n4404 net3271 VDD pmos w=2u l=1u
M10912 net3271 n4403 VDD VDD pmos w=2u l=1u
M10913 n4404 net3272 VSS VSS nmos w=1u l=1u
M10914 net3273 n4346 VSS VSS nmos w=1u l=1u
M10915 net3272 n4347 net3273 VSS nmos w=1u l=1u
M10916 net3272 n4346 VDD VDD pmos w=2u l=1u
M10917 net3272 n4347 VDD VDD pmos w=2u l=1u
M10918 n4404 net3272 VDD VDD pmos w=2u l=1u
M10919 n4403 n4345 VDD VDD pmos w=2u l=1u
M10920 n4403 n4345 VSS VSS nmos w=1u l=1u
M10921 n4339 n4406 VSS VSS nmos w=1u l=1u
M10922 n4339 n4405 VSS VSS nmos w=1u l=1u
M10923 n4339 n4406 net3274 VDD pmos w=2u l=1u
M10924 net3274 n4405 VDD VDD pmos w=2u l=1u
M10925 n4406 n4408 VSS VSS nmos w=1u l=1u
M10926 n4406 n4407 VSS VSS nmos w=1u l=1u
M10927 n4406 n4408 net3275 VDD pmos w=2u l=1u
M10928 net3275 n4407 VDD VDD pmos w=2u l=1u
M10929 n4407 n4337 VDD VDD pmos w=2u l=1u
M10930 n4407 n4337 VSS VSS nmos w=1u l=1u
M10931 n4405 n4335 VDD VDD pmos w=2u l=1u
M10932 n4405 n4335 VSS VSS nmos w=1u l=1u
M10933 n4329 n4410 VSS VSS nmos w=1u l=1u
M10934 n4329 n4409 VSS VSS nmos w=1u l=1u
M10935 n4329 n4410 net3276 VDD pmos w=2u l=1u
M10936 net3276 n4409 VDD VDD pmos w=2u l=1u
M10937 n4410 n4412 VSS VSS nmos w=1u l=1u
M10938 n4410 n4411 VSS VSS nmos w=1u l=1u
M10939 n4410 n4412 net3277 VDD pmos w=2u l=1u
M10940 net3277 n4411 VDD VDD pmos w=2u l=1u
M10941 n4411 n4328 VDD VDD pmos w=2u l=1u
M10942 n4411 n4328 VSS VSS nmos w=1u l=1u
M10943 n4409 n4326 VDD VDD pmos w=2u l=1u
M10944 n4409 n4326 VSS VSS nmos w=1u l=1u
M10945 n4320 n4414 VSS VSS nmos w=1u l=1u
M10946 n4320 n4413 VSS VSS nmos w=1u l=1u
M10947 n4320 n4414 net3278 VDD pmos w=2u l=1u
M10948 net3278 n4413 VDD VDD pmos w=2u l=1u
M10949 n4414 n4318 VSS VSS nmos w=1u l=1u
M10950 n4414 n4319 VSS VSS nmos w=1u l=1u
M10951 n4414 n4318 net3279 VDD pmos w=2u l=1u
M10952 net3279 n4319 VDD VDD pmos w=2u l=1u
M10953 n4413 n4317 VDD VDD pmos w=2u l=1u
M10954 n4413 n4317 VSS VSS nmos w=1u l=1u
M10955 net3280 n4319 VSS VSS nmos w=1u l=1u
M10956 net3281 n4415 VSS VSS nmos w=1u l=1u
M10957 N4241 net3282 VSS VSS nmos w=1u l=1u
M10958 net3282 n4319 net3283 VSS nmos w=1u l=1u
M10959 net3282 net3280 net3281 VSS nmos w=1u l=1u
M10960 net3283 net3281 VSS VSS nmos w=1u l=1u
M10961 net3282 net3280 net3284 VDD pmos w=2u l=1u
M10962 net3280 n4319 VDD VDD pmos w=2u l=1u
M10963 net3281 n4319 net3282 VDD pmos w=2u l=1u
M10964 net3281 n4415 VDD VDD pmos w=2u l=1u
M10965 N4241 net3282 VDD VDD pmos w=2u l=1u
M10966 net3284 net3281 VDD VDD pmos w=2u l=1u
M10967 n4319 n2525 VSS VSS nmos w=1u l=1u
M10968 n4319 n3929 VSS VSS nmos w=1u l=1u
M10969 n4319 n2525 net3285 VDD pmos w=2u l=1u
M10970 net3285 n3929 VDD VDD pmos w=2u l=1u
M10971 n2525 N426 VDD VDD pmos w=2u l=1u
M10972 n2525 N426 VSS VSS nmos w=1u l=1u
M10973 n4415 n4318 VDD VDD pmos w=2u l=1u
M10974 n4415 n4318 VSS VSS nmos w=1u l=1u
M10975 n4318 n4317 net3286 VSS nmos w=1u l=1u
M10976 net3286 n4416 VSS VSS nmos w=1u l=1u
M10977 n4318 n4317 VDD VDD pmos w=2u l=1u
M10978 n4318 n4416 VDD VDD pmos w=2u l=1u
M10979 n4317 n4418 net3287 VSS nmos w=1u l=1u
M10980 net3287 n4417 VSS VSS nmos w=1u l=1u
M10981 n4317 n4418 VDD VDD pmos w=2u l=1u
M10982 n4317 n4417 VDD VDD pmos w=2u l=1u
M10983 n4418 n4420 net3288 VSS nmos w=1u l=1u
M10984 net3288 n4419 VSS VSS nmos w=1u l=1u
M10985 n4418 n4420 VDD VDD pmos w=2u l=1u
M10986 n4418 n4419 VDD VDD pmos w=2u l=1u
M10987 n4419 net3289 VSS VSS nmos w=1u l=1u
M10988 net3289 n4421 VSS VSS nmos w=1u l=1u
M10989 net3289 n4422 VSS VSS nmos w=1u l=1u
M10990 net3289 n4422 net3290 VDD pmos w=2u l=1u
M10991 n4419 net3289 VDD VDD pmos w=2u l=1u
M10992 net3290 n4421 VDD VDD pmos w=2u l=1u
M10993 net3291 n4327 VSS VSS nmos w=1u l=1u
M10994 net3292 n4328 VSS VSS nmos w=1u l=1u
M10995 n4417 net3293 VSS VSS nmos w=1u l=1u
M10996 net3293 n4327 net3294 VSS nmos w=1u l=1u
M10997 net3293 net3291 net3292 VSS nmos w=1u l=1u
M10998 net3294 net3292 VSS VSS nmos w=1u l=1u
M10999 net3293 net3291 net3295 VDD pmos w=2u l=1u
M11000 net3291 n4327 VDD VDD pmos w=2u l=1u
M11001 net3292 n4327 net3293 VDD pmos w=2u l=1u
M11002 net3292 n4328 VDD VDD pmos w=2u l=1u
M11003 n4417 net3293 VDD VDD pmos w=2u l=1u
M11004 net3295 net3292 VDD VDD pmos w=2u l=1u
M11005 n4327 n4412 VDD VDD pmos w=2u l=1u
M11006 n4327 n4412 VSS VSS nmos w=1u l=1u
M11007 n4416 n4424 net3296 VSS nmos w=1u l=1u
M11008 net3296 n4423 VSS VSS nmos w=1u l=1u
M11009 n4416 n4424 VDD VDD pmos w=2u l=1u
M11010 n4416 n4423 VDD VDD pmos w=2u l=1u
M11011 net3297 n4328 VSS VSS nmos w=1u l=1u
M11012 net3298 n4412 VSS VSS nmos w=1u l=1u
M11013 n4424 net3299 VSS VSS nmos w=1u l=1u
M11014 net3299 n4328 net3300 VSS nmos w=1u l=1u
M11015 net3299 net3297 net3298 VSS nmos w=1u l=1u
M11016 net3300 net3298 VSS VSS nmos w=1u l=1u
M11017 net3299 net3297 net3301 VDD pmos w=2u l=1u
M11018 net3297 n4328 VDD VDD pmos w=2u l=1u
M11019 net3298 n4328 net3299 VDD pmos w=2u l=1u
M11020 net3298 n4412 VDD VDD pmos w=2u l=1u
M11021 n4424 net3299 VDD VDD pmos w=2u l=1u
M11022 net3301 net3298 VDD VDD pmos w=2u l=1u
M11023 n4328 N409 net3302 VSS nmos w=1u l=1u
M11024 net3302 N18 VSS VSS nmos w=1u l=1u
M11025 n4328 N409 VDD VDD pmos w=2u l=1u
M11026 n4328 N18 VDD VDD pmos w=2u l=1u
M11027 n4412 n4326 net3303 VSS nmos w=1u l=1u
M11028 net3303 n4425 VSS VSS nmos w=1u l=1u
M11029 n4412 n4326 VDD VDD pmos w=2u l=1u
M11030 n4412 n4425 VDD VDD pmos w=2u l=1u
M11031 n4326 n4427 net3304 VSS nmos w=1u l=1u
M11032 net3304 n4426 VSS VSS nmos w=1u l=1u
M11033 n4326 n4427 VDD VDD pmos w=2u l=1u
M11034 n4326 n4426 VDD VDD pmos w=2u l=1u
M11035 n4427 n4429 net3305 VSS nmos w=1u l=1u
M11036 net3305 n4428 VSS VSS nmos w=1u l=1u
M11037 n4427 n4429 VDD VDD pmos w=2u l=1u
M11038 n4427 n4428 VDD VDD pmos w=2u l=1u
M11039 n4428 n4431 net3306 VSS nmos w=1u l=1u
M11040 net3306 n4430 VSS VSS nmos w=1u l=1u
M11041 n4428 n4431 VDD VDD pmos w=2u l=1u
M11042 n4428 n4430 VDD VDD pmos w=2u l=1u
M11043 net3307 n4336 VSS VSS nmos w=1u l=1u
M11044 net3308 n4337 VSS VSS nmos w=1u l=1u
M11045 n4426 net3309 VSS VSS nmos w=1u l=1u
M11046 net3309 n4336 net3310 VSS nmos w=1u l=1u
M11047 net3309 net3307 net3308 VSS nmos w=1u l=1u
M11048 net3310 net3308 VSS VSS nmos w=1u l=1u
M11049 net3309 net3307 net3311 VDD pmos w=2u l=1u
M11050 net3307 n4336 VDD VDD pmos w=2u l=1u
M11051 net3308 n4336 net3309 VDD pmos w=2u l=1u
M11052 net3308 n4337 VDD VDD pmos w=2u l=1u
M11053 n4426 net3309 VDD VDD pmos w=2u l=1u
M11054 net3311 net3308 VDD VDD pmos w=2u l=1u
M11055 n4336 n4408 VDD VDD pmos w=2u l=1u
M11056 n4336 n4408 VSS VSS nmos w=1u l=1u
M11057 n4425 n4433 net3312 VSS nmos w=1u l=1u
M11058 net3312 n4432 VSS VSS nmos w=1u l=1u
M11059 n4425 n4433 VDD VDD pmos w=2u l=1u
M11060 n4425 n4432 VDD VDD pmos w=2u l=1u
M11061 net3313 n4337 VSS VSS nmos w=1u l=1u
M11062 net3314 n4408 VSS VSS nmos w=1u l=1u
M11063 n4433 net3315 VSS VSS nmos w=1u l=1u
M11064 net3315 n4337 net3316 VSS nmos w=1u l=1u
M11065 net3315 net3313 net3314 VSS nmos w=1u l=1u
M11066 net3316 net3314 VSS VSS nmos w=1u l=1u
M11067 net3315 net3313 net3317 VDD pmos w=2u l=1u
M11068 net3313 n4337 VDD VDD pmos w=2u l=1u
M11069 net3314 n4337 net3315 VDD pmos w=2u l=1u
M11070 net3314 n4408 VDD VDD pmos w=2u l=1u
M11071 n4433 net3315 VDD VDD pmos w=2u l=1u
M11072 net3317 net3314 VDD VDD pmos w=2u l=1u
M11073 n4337 N392 net3318 VSS nmos w=1u l=1u
M11074 net3318 N35 VSS VSS nmos w=1u l=1u
M11075 n4337 N392 VDD VDD pmos w=2u l=1u
M11076 n4337 N35 VDD VDD pmos w=2u l=1u
M11077 n4408 n4335 net3319 VSS nmos w=1u l=1u
M11078 net3319 n4434 VSS VSS nmos w=1u l=1u
M11079 n4408 n4335 VDD VDD pmos w=2u l=1u
M11080 n4408 n4434 VDD VDD pmos w=2u l=1u
M11081 n4335 n4436 net3320 VSS nmos w=1u l=1u
M11082 net3320 n4435 VSS VSS nmos w=1u l=1u
M11083 n4335 n4436 VDD VDD pmos w=2u l=1u
M11084 n4335 n4435 VDD VDD pmos w=2u l=1u
M11085 n4436 n4438 net3321 VSS nmos w=1u l=1u
M11086 net3321 n4437 VSS VSS nmos w=1u l=1u
M11087 n4436 n4438 VDD VDD pmos w=2u l=1u
M11088 n4436 n4437 VDD VDD pmos w=2u l=1u
M11089 n4437 n4440 net3322 VSS nmos w=1u l=1u
M11090 net3322 n4439 VSS VSS nmos w=1u l=1u
M11091 n4437 n4440 VDD VDD pmos w=2u l=1u
M11092 n4437 n4439 VDD VDD pmos w=2u l=1u
M11093 net3323 n4346 VSS VSS nmos w=1u l=1u
M11094 net3324 n4347 VSS VSS nmos w=1u l=1u
M11095 n4435 net3325 VSS VSS nmos w=1u l=1u
M11096 net3325 n4346 net3326 VSS nmos w=1u l=1u
M11097 net3325 net3323 net3324 VSS nmos w=1u l=1u
M11098 net3326 net3324 VSS VSS nmos w=1u l=1u
M11099 net3325 net3323 net3327 VDD pmos w=2u l=1u
M11100 net3323 n4346 VDD VDD pmos w=2u l=1u
M11101 net3324 n4346 net3325 VDD pmos w=2u l=1u
M11102 net3324 n4347 VDD VDD pmos w=2u l=1u
M11103 n4435 net3325 VDD VDD pmos w=2u l=1u
M11104 net3327 net3324 VDD VDD pmos w=2u l=1u
M11105 n4346 n4441 VDD VDD pmos w=2u l=1u
M11106 n4346 n4441 VSS VSS nmos w=1u l=1u
M11107 n4434 n4443 net3328 VSS nmos w=1u l=1u
M11108 net3328 n4442 VSS VSS nmos w=1u l=1u
M11109 n4434 n4443 VDD VDD pmos w=2u l=1u
M11110 n4434 n4442 VDD VDD pmos w=2u l=1u
M11111 net3329 n4347 VSS VSS nmos w=1u l=1u
M11112 net3330 n4441 VSS VSS nmos w=1u l=1u
M11113 n4443 net3331 VSS VSS nmos w=1u l=1u
M11114 net3331 n4347 net3332 VSS nmos w=1u l=1u
M11115 net3331 net3329 net3330 VSS nmos w=1u l=1u
M11116 net3332 net3330 VSS VSS nmos w=1u l=1u
M11117 net3331 net3329 net3333 VDD pmos w=2u l=1u
M11118 net3329 n4347 VDD VDD pmos w=2u l=1u
M11119 net3330 n4347 net3331 VDD pmos w=2u l=1u
M11120 net3330 n4441 VDD VDD pmos w=2u l=1u
M11121 n4443 net3331 VDD VDD pmos w=2u l=1u
M11122 net3333 net3330 VDD VDD pmos w=2u l=1u
M11123 n4347 N375 net3334 VSS nmos w=1u l=1u
M11124 net3334 N52 VSS VSS nmos w=1u l=1u
M11125 n4347 N375 VDD VDD pmos w=2u l=1u
M11126 n4347 N52 VDD VDD pmos w=2u l=1u
M11127 n4441 n4345 net3335 VSS nmos w=1u l=1u
M11128 net3335 n4444 VSS VSS nmos w=1u l=1u
M11129 n4441 n4345 VDD VDD pmos w=2u l=1u
M11130 n4441 n4444 VDD VDD pmos w=2u l=1u
M11131 n4345 n4446 net3336 VSS nmos w=1u l=1u
M11132 net3336 n4445 VSS VSS nmos w=1u l=1u
M11133 n4345 n4446 VDD VDD pmos w=2u l=1u
M11134 n4345 n4445 VDD VDD pmos w=2u l=1u
M11135 n4446 n4448 net3337 VSS nmos w=1u l=1u
M11136 net3337 n4447 VSS VSS nmos w=1u l=1u
M11137 n4446 n4448 VDD VDD pmos w=2u l=1u
M11138 n4446 n4447 VDD VDD pmos w=2u l=1u
M11139 n4447 net3338 VSS VSS nmos w=1u l=1u
M11140 net3338 n4449 VSS VSS nmos w=1u l=1u
M11141 net3338 n4450 VSS VSS nmos w=1u l=1u
M11142 net3338 n4450 net3339 VDD pmos w=2u l=1u
M11143 n4447 net3338 VDD VDD pmos w=2u l=1u
M11144 net3339 n4449 VDD VDD pmos w=2u l=1u
M11145 net3340 n4356 VSS VSS nmos w=1u l=1u
M11146 net3341 n4357 VSS VSS nmos w=1u l=1u
M11147 n4445 net3342 VSS VSS nmos w=1u l=1u
M11148 net3342 n4356 net3343 VSS nmos w=1u l=1u
M11149 net3342 net3340 net3341 VSS nmos w=1u l=1u
M11150 net3343 net3341 VSS VSS nmos w=1u l=1u
M11151 net3342 net3340 net3344 VDD pmos w=2u l=1u
M11152 net3340 n4356 VDD VDD pmos w=2u l=1u
M11153 net3341 n4356 net3342 VDD pmos w=2u l=1u
M11154 net3341 n4357 VDD VDD pmos w=2u l=1u
M11155 n4445 net3342 VDD VDD pmos w=2u l=1u
M11156 net3344 net3341 VDD VDD pmos w=2u l=1u
M11157 n4357 n4451 VDD VDD pmos w=2u l=1u
M11158 n4357 n4451 VSS VSS nmos w=1u l=1u
M11159 n4444 n4453 net3345 VSS nmos w=1u l=1u
M11160 net3345 n4452 VSS VSS nmos w=1u l=1u
M11161 n4444 n4453 VDD VDD pmos w=2u l=1u
M11162 n4444 n4452 VDD VDD pmos w=2u l=1u
M11163 net3346 n4451 VSS VSS nmos w=1u l=1u
M11164 net3347 n4356 VSS VSS nmos w=1u l=1u
M11165 n4453 net3348 VSS VSS nmos w=1u l=1u
M11166 net3348 n4451 net3349 VSS nmos w=1u l=1u
M11167 net3348 net3346 net3347 VSS nmos w=1u l=1u
M11168 net3349 net3347 VSS VSS nmos w=1u l=1u
M11169 net3348 net3346 net3350 VDD pmos w=2u l=1u
M11170 net3346 n4451 VDD VDD pmos w=2u l=1u
M11171 net3347 n4451 net3348 VDD pmos w=2u l=1u
M11172 net3347 n4356 VDD VDD pmos w=2u l=1u
M11173 n4453 net3348 VDD VDD pmos w=2u l=1u
M11174 net3350 net3347 VDD VDD pmos w=2u l=1u
M11175 n4451 N358 net3351 VSS nmos w=1u l=1u
M11176 net3351 N69 VSS VSS nmos w=1u l=1u
M11177 n4451 N358 VDD VDD pmos w=2u l=1u
M11178 n4451 N69 VDD VDD pmos w=2u l=1u
M11179 n4356 n4355 net3352 VSS nmos w=1u l=1u
M11180 net3352 n4454 VSS VSS nmos w=1u l=1u
M11181 n4356 n4355 VDD VDD pmos w=2u l=1u
M11182 n4356 n4454 VDD VDD pmos w=2u l=1u
M11183 n4355 n4456 net3353 VSS nmos w=1u l=1u
M11184 net3353 n4455 VSS VSS nmos w=1u l=1u
M11185 n4355 n4456 VDD VDD pmos w=2u l=1u
M11186 n4355 n4455 VDD VDD pmos w=2u l=1u
M11187 n4456 n4458 net3354 VSS nmos w=1u l=1u
M11188 net3354 n4457 VSS VSS nmos w=1u l=1u
M11189 n4456 n4458 VDD VDD pmos w=2u l=1u
M11190 n4456 n4457 VDD VDD pmos w=2u l=1u
M11191 n4457 n4460 net3355 VSS nmos w=1u l=1u
M11192 net3355 n4459 VSS VSS nmos w=1u l=1u
M11193 n4457 n4460 VDD VDD pmos w=2u l=1u
M11194 n4457 n4459 VDD VDD pmos w=2u l=1u
M11195 net3356 n4366 VSS VSS nmos w=1u l=1u
M11196 net3357 n4367 VSS VSS nmos w=1u l=1u
M11197 n4455 net3358 VSS VSS nmos w=1u l=1u
M11198 net3358 n4366 net3359 VSS nmos w=1u l=1u
M11199 net3358 net3356 net3357 VSS nmos w=1u l=1u
M11200 net3359 net3357 VSS VSS nmos w=1u l=1u
M11201 net3358 net3356 net3360 VDD pmos w=2u l=1u
M11202 net3356 n4366 VDD VDD pmos w=2u l=1u
M11203 net3357 n4366 net3358 VDD pmos w=2u l=1u
M11204 net3357 n4367 VDD VDD pmos w=2u l=1u
M11205 n4455 net3358 VDD VDD pmos w=2u l=1u
M11206 net3360 net3357 VDD VDD pmos w=2u l=1u
M11207 n4366 n4461 VDD VDD pmos w=2u l=1u
M11208 n4366 n4461 VSS VSS nmos w=1u l=1u
M11209 n4454 n4463 net3361 VSS nmos w=1u l=1u
M11210 net3361 n4462 VSS VSS nmos w=1u l=1u
M11211 n4454 n4463 VDD VDD pmos w=2u l=1u
M11212 n4454 n4462 VDD VDD pmos w=2u l=1u
M11213 net3362 n4367 VSS VSS nmos w=1u l=1u
M11214 net3363 n4461 VSS VSS nmos w=1u l=1u
M11215 n4463 net3364 VSS VSS nmos w=1u l=1u
M11216 net3364 n4367 net3365 VSS nmos w=1u l=1u
M11217 net3364 net3362 net3363 VSS nmos w=1u l=1u
M11218 net3365 net3363 VSS VSS nmos w=1u l=1u
M11219 net3364 net3362 net3366 VDD pmos w=2u l=1u
M11220 net3362 n4367 VDD VDD pmos w=2u l=1u
M11221 net3363 n4367 net3364 VDD pmos w=2u l=1u
M11222 net3363 n4461 VDD VDD pmos w=2u l=1u
M11223 n4463 net3364 VDD VDD pmos w=2u l=1u
M11224 net3366 net3363 VDD VDD pmos w=2u l=1u
M11225 n4367 N341 net3367 VSS nmos w=1u l=1u
M11226 net3367 N86 VSS VSS nmos w=1u l=1u
M11227 n4367 N341 VDD VDD pmos w=2u l=1u
M11228 n4367 N86 VDD VDD pmos w=2u l=1u
M11229 n4461 n4365 net3368 VSS nmos w=1u l=1u
M11230 net3368 n4464 VSS VSS nmos w=1u l=1u
M11231 n4461 n4365 VDD VDD pmos w=2u l=1u
M11232 n4461 n4464 VDD VDD pmos w=2u l=1u
M11233 n4365 n4466 net3369 VSS nmos w=1u l=1u
M11234 net3369 n4465 VSS VSS nmos w=1u l=1u
M11235 n4365 n4466 VDD VDD pmos w=2u l=1u
M11236 n4365 n4465 VDD VDD pmos w=2u l=1u
M11237 n4466 net3370 VSS VSS nmos w=1u l=1u
M11238 net3370 n4467 VSS VSS nmos w=1u l=1u
M11239 net3370 n4468 VSS VSS nmos w=1u l=1u
M11240 net3370 n4468 net3371 VDD pmos w=2u l=1u
M11241 n4466 net3370 VDD VDD pmos w=2u l=1u
M11242 net3371 n4467 VDD VDD pmos w=2u l=1u
M11243 n4465 net3372 VSS VSS nmos w=1u l=1u
M11244 net3373 n4469 VSS VSS nmos w=1u l=1u
M11245 net3372 n4398 net3373 VSS nmos w=1u l=1u
M11246 net3372 n4469 VDD VDD pmos w=2u l=1u
M11247 net3372 n4398 VDD VDD pmos w=2u l=1u
M11248 n4465 net3372 VDD VDD pmos w=2u l=1u
M11249 n4464 n4471 net3374 VSS nmos w=1u l=1u
M11250 net3374 n4470 VSS VSS nmos w=1u l=1u
M11251 n4464 n4471 VDD VDD pmos w=2u l=1u
M11252 n4464 n4470 VDD VDD pmos w=2u l=1u
M11253 n4471 n4398 net3375 VSS nmos w=1u l=1u
M11254 net3375 n4469 VSS VSS nmos w=1u l=1u
M11255 n4471 n4398 VDD VDD pmos w=2u l=1u
M11256 n4471 n4469 VDD VDD pmos w=2u l=1u
M11257 n4398 n4473 net3376 VSS nmos w=1u l=1u
M11258 net3376 n4472 VSS VSS nmos w=1u l=1u
M11259 n4398 n4473 VDD VDD pmos w=2u l=1u
M11260 n4398 n4472 VDD VDD pmos w=2u l=1u
M11261 n4473 N324 net3377 VSS nmos w=1u l=1u
M11262 net3377 N103 VSS VSS nmos w=1u l=1u
M11263 n4473 N324 VDD VDD pmos w=2u l=1u
M11264 n4473 N103 VDD VDD pmos w=2u l=1u
M11265 n4469 N103 net3378 VSS nmos w=1u l=1u
M11266 net3378 n4474 VSS VSS nmos w=1u l=1u
M11267 n4469 N103 VDD VDD pmos w=2u l=1u
M11268 n4469 n4474 VDD VDD pmos w=2u l=1u
M11269 n4474 n3257 VSS VSS nmos w=1u l=1u
M11270 n4474 n4472 VSS VSS nmos w=1u l=1u
M11271 n4474 n3257 net3379 VDD pmos w=2u l=1u
M11272 net3379 n4472 VDD VDD pmos w=2u l=1u
M11273 n4472 n4375 VSS VSS nmos w=1u l=1u
M11274 n4472 n4475 VSS VSS nmos w=1u l=1u
M11275 n4472 n4375 net3380 VDD pmos w=2u l=1u
M11276 net3380 n4475 VDD VDD pmos w=2u l=1u
M11277 n4375 n4477 VSS VSS nmos w=1u l=1u
M11278 n4375 n4476 VSS VSS nmos w=1u l=1u
M11279 n4375 n4477 net3381 VDD pmos w=2u l=1u
M11280 net3381 n4476 VDD VDD pmos w=2u l=1u
M11281 n4475 net3382 VSS VSS nmos w=1u l=1u
M11282 net3383 n4476 VSS VSS nmos w=1u l=1u
M11283 net3382 n4477 net3383 VSS nmos w=1u l=1u
M11284 net3382 n4476 VDD VDD pmos w=2u l=1u
M11285 net3382 n4477 VDD VDD pmos w=2u l=1u
M11286 n4475 net3382 VDD VDD pmos w=2u l=1u
M11287 n4476 n4478 net3384 VSS nmos w=1u l=1u
M11288 net3384 n4396 VSS VSS nmos w=1u l=1u
M11289 n4476 n4478 VDD VDD pmos w=2u l=1u
M11290 n4476 n4396 VDD VDD pmos w=2u l=1u
M11291 n4478 N120 net3385 VSS nmos w=1u l=1u
M11292 net3385 n4479 VSS VSS nmos w=1u l=1u
M11293 n4478 N120 VDD VDD pmos w=2u l=1u
M11294 n4478 n4479 VDD VDD pmos w=2u l=1u
M11295 n4479 n3411 VSS VSS nmos w=1u l=1u
M11296 n4479 n4480 VSS VSS nmos w=1u l=1u
M11297 n4479 n3411 net3386 VDD pmos w=2u l=1u
M11298 net3386 n4480 VDD VDD pmos w=2u l=1u
M11299 n4396 n4481 net3387 VSS nmos w=1u l=1u
M11300 net3387 n4480 VSS VSS nmos w=1u l=1u
M11301 n4396 n4481 VDD VDD pmos w=2u l=1u
M11302 n4396 n4480 VDD VDD pmos w=2u l=1u
M11303 n4481 N307 net3388 VSS nmos w=1u l=1u
M11304 net3388 N120 VSS VSS nmos w=1u l=1u
M11305 n4481 N307 VDD VDD pmos w=2u l=1u
M11306 n4481 N120 VDD VDD pmos w=2u l=1u
M11307 n4480 net3389 VSS VSS nmos w=1u l=1u
M11308 net3390 n4482 VSS VSS nmos w=1u l=1u
M11309 net3389 n4397 net3390 VSS nmos w=1u l=1u
M11310 net3389 n4482 VDD VDD pmos w=2u l=1u
M11311 net3389 n4397 VDD VDD pmos w=2u l=1u
M11312 n4480 net3389 VDD VDD pmos w=2u l=1u
M11313 n4482 n4390 net3391 VSS nmos w=1u l=1u
M11314 net3391 n4483 VSS VSS nmos w=1u l=1u
M11315 n4482 n4390 VDD VDD pmos w=2u l=1u
M11316 n4482 n4483 VDD VDD pmos w=2u l=1u
M11317 n4397 n4485 net3392 VSS nmos w=1u l=1u
M11318 net3392 n4484 VSS VSS nmos w=1u l=1u
M11319 n4397 n4485 VDD VDD pmos w=2u l=1u
M11320 n4397 n4484 VDD VDD pmos w=2u l=1u
M11321 n4485 n4390 net3393 VSS nmos w=1u l=1u
M11322 net3393 n4486 VSS VSS nmos w=1u l=1u
M11323 n4485 n4390 VDD VDD pmos w=2u l=1u
M11324 n4485 n4486 VDD VDD pmos w=2u l=1u
M11325 n4390 N154 net3394 VSS nmos w=1u l=1u
M11326 net3394 n4487 VSS VSS nmos w=1u l=1u
M11327 n4390 N154 VDD VDD pmos w=2u l=1u
M11328 n4390 n4487 VDD VDD pmos w=2u l=1u
M11329 n4487 net3395 VSS VSS nmos w=1u l=1u
M11330 net3396 N137 VSS VSS nmos w=1u l=1u
M11331 net3395 n3741 net3396 VSS nmos w=1u l=1u
M11332 net3395 N137 VDD VDD pmos w=2u l=1u
M11333 net3395 n3741 VDD VDD pmos w=2u l=1u
M11334 n4487 net3395 VDD VDD pmos w=2u l=1u
M11335 n4486 n4489 net3397 VSS nmos w=1u l=1u
M11336 net3397 n4488 VSS VSS nmos w=1u l=1u
M11337 n4486 n4489 VDD VDD pmos w=2u l=1u
M11338 n4486 n4488 VDD VDD pmos w=2u l=1u
M11339 n4489 N273 net3398 VSS nmos w=1u l=1u
M11340 net3398 N154 VSS VSS nmos w=1u l=1u
M11341 n4489 N273 VDD VDD pmos w=2u l=1u
M11342 n4489 N154 VDD VDD pmos w=2u l=1u
M11343 n4488 N290 net3399 VSS nmos w=1u l=1u
M11344 net3399 N137 VSS VSS nmos w=1u l=1u
M11345 n4488 N290 VDD VDD pmos w=2u l=1u
M11346 n4488 N137 VDD VDD pmos w=2u l=1u
M11347 n4477 net3400 VSS VSS nmos w=1u l=1u
M11348 net3401 n4491 VSS VSS nmos w=1u l=1u
M11349 net3400 n4490 net3401 VSS nmos w=1u l=1u
M11350 net3400 n4491 VDD VDD pmos w=2u l=1u
M11351 net3400 n4490 VDD VDD pmos w=2u l=1u
M11352 n4477 net3400 VDD VDD pmos w=2u l=1u
M11353 n4470 n4467 VSS VSS nmos w=1u l=1u
M11354 n4470 n4468 VSS VSS nmos w=1u l=1u
M11355 n4470 n4467 net3402 VDD pmos w=2u l=1u
M11356 net3402 n4468 VDD VDD pmos w=2u l=1u
M11357 n4467 n4492 VDD VDD pmos w=2u l=1u
M11358 n4467 n4492 VSS VSS nmos w=1u l=1u
M11359 n4462 n4494 VSS VSS nmos w=1u l=1u
M11360 n4462 n4493 VSS VSS nmos w=1u l=1u
M11361 n4462 n4494 net3403 VDD pmos w=2u l=1u
M11362 net3403 n4493 VDD VDD pmos w=2u l=1u
M11363 n4494 net3404 VSS VSS nmos w=1u l=1u
M11364 net3405 n4459 VSS VSS nmos w=1u l=1u
M11365 net3404 n4460 net3405 VSS nmos w=1u l=1u
M11366 net3404 n4459 VDD VDD pmos w=2u l=1u
M11367 net3404 n4460 VDD VDD pmos w=2u l=1u
M11368 n4494 net3404 VDD VDD pmos w=2u l=1u
M11369 n4493 n4458 VDD VDD pmos w=2u l=1u
M11370 n4493 n4458 VSS VSS nmos w=1u l=1u
M11371 n4452 n4496 VSS VSS nmos w=1u l=1u
M11372 n4452 n4495 VSS VSS nmos w=1u l=1u
M11373 n4452 n4496 net3406 VDD pmos w=2u l=1u
M11374 net3406 n4495 VDD VDD pmos w=2u l=1u
M11375 n4496 n4449 VSS VSS nmos w=1u l=1u
M11376 n4496 n4450 VSS VSS nmos w=1u l=1u
M11377 n4496 n4449 net3407 VDD pmos w=2u l=1u
M11378 net3407 n4450 VDD VDD pmos w=2u l=1u
M11379 n4495 n4448 VDD VDD pmos w=2u l=1u
M11380 n4495 n4448 VSS VSS nmos w=1u l=1u
M11381 n4442 n4498 VSS VSS nmos w=1u l=1u
M11382 n4442 n4497 VSS VSS nmos w=1u l=1u
M11383 n4442 n4498 net3408 VDD pmos w=2u l=1u
M11384 net3408 n4497 VDD VDD pmos w=2u l=1u
M11385 n4498 n4500 VSS VSS nmos w=1u l=1u
M11386 n4498 n4499 VSS VSS nmos w=1u l=1u
M11387 n4498 n4500 net3409 VDD pmos w=2u l=1u
M11388 net3409 n4499 VDD VDD pmos w=2u l=1u
M11389 n4499 n4440 VDD VDD pmos w=2u l=1u
M11390 n4499 n4440 VSS VSS nmos w=1u l=1u
M11391 n4497 n4438 VDD VDD pmos w=2u l=1u
M11392 n4497 n4438 VSS VSS nmos w=1u l=1u
M11393 n4432 n4502 VSS VSS nmos w=1u l=1u
M11394 n4432 n4501 VSS VSS nmos w=1u l=1u
M11395 n4432 n4502 net3410 VDD pmos w=2u l=1u
M11396 net3410 n4501 VDD VDD pmos w=2u l=1u
M11397 n4502 n4504 VSS VSS nmos w=1u l=1u
M11398 n4502 n4503 VSS VSS nmos w=1u l=1u
M11399 n4502 n4504 net3411 VDD pmos w=2u l=1u
M11400 net3411 n4503 VDD VDD pmos w=2u l=1u
M11401 n4503 n4431 VDD VDD pmos w=2u l=1u
M11402 n4503 n4431 VSS VSS nmos w=1u l=1u
M11403 n4501 n4429 VDD VDD pmos w=2u l=1u
M11404 n4501 n4429 VSS VSS nmos w=1u l=1u
M11405 n4423 n4506 VSS VSS nmos w=1u l=1u
M11406 n4423 n4505 VSS VSS nmos w=1u l=1u
M11407 n4423 n4506 net3412 VDD pmos w=2u l=1u
M11408 net3412 n4505 VDD VDD pmos w=2u l=1u
M11409 n4506 n4421 VSS VSS nmos w=1u l=1u
M11410 n4506 n4422 VSS VSS nmos w=1u l=1u
M11411 n4506 n4421 net3413 VDD pmos w=2u l=1u
M11412 net3413 n4422 VDD VDD pmos w=2u l=1u
M11413 n4505 n4420 VDD VDD pmos w=2u l=1u
M11414 n4505 n4420 VSS VSS nmos w=1u l=1u
M11415 net3414 n4422 VSS VSS nmos w=1u l=1u
M11416 net3415 n4507 VSS VSS nmos w=1u l=1u
M11417 N3895 net3416 VSS VSS nmos w=1u l=1u
M11418 net3416 n4422 net3417 VSS nmos w=1u l=1u
M11419 net3416 net3414 net3415 VSS nmos w=1u l=1u
M11420 net3417 net3415 VSS VSS nmos w=1u l=1u
M11421 net3416 net3414 net3418 VDD pmos w=2u l=1u
M11422 net3414 n4422 VDD VDD pmos w=2u l=1u
M11423 net3415 n4422 net3416 VDD pmos w=2u l=1u
M11424 net3415 n4507 VDD VDD pmos w=2u l=1u
M11425 N3895 net3416 VDD VDD pmos w=2u l=1u
M11426 net3418 net3415 VDD VDD pmos w=2u l=1u
M11427 n4422 n2617 VSS VSS nmos w=1u l=1u
M11428 n4422 n3929 VSS VSS nmos w=1u l=1u
M11429 n4422 n2617 net3419 VDD pmos w=2u l=1u
M11430 net3419 n3929 VDD VDD pmos w=2u l=1u
M11431 n2617 N409 VDD VDD pmos w=2u l=1u
M11432 n2617 N409 VSS VSS nmos w=1u l=1u
M11433 n4507 n4421 VDD VDD pmos w=2u l=1u
M11434 n4507 n4421 VSS VSS nmos w=1u l=1u
M11435 n4421 n4420 net3420 VSS nmos w=1u l=1u
M11436 net3420 n4508 VSS VSS nmos w=1u l=1u
M11437 n4421 n4420 VDD VDD pmos w=2u l=1u
M11438 n4421 n4508 VDD VDD pmos w=2u l=1u
M11439 n4420 n4510 net3421 VSS nmos w=1u l=1u
M11440 net3421 n4509 VSS VSS nmos w=1u l=1u
M11441 n4420 n4510 VDD VDD pmos w=2u l=1u
M11442 n4420 n4509 VDD VDD pmos w=2u l=1u
M11443 n4510 n4512 net3422 VSS nmos w=1u l=1u
M11444 net3422 n4511 VSS VSS nmos w=1u l=1u
M11445 n4510 n4512 VDD VDD pmos w=2u l=1u
M11446 n4510 n4511 VDD VDD pmos w=2u l=1u
M11447 n4511 net3423 VSS VSS nmos w=1u l=1u
M11448 net3423 n4513 VSS VSS nmos w=1u l=1u
M11449 net3423 n4514 VSS VSS nmos w=1u l=1u
M11450 net3423 n4514 net3424 VDD pmos w=2u l=1u
M11451 n4511 net3423 VDD VDD pmos w=2u l=1u
M11452 net3424 n4513 VDD VDD pmos w=2u l=1u
M11453 net3425 n4430 VSS VSS nmos w=1u l=1u
M11454 net3426 n4431 VSS VSS nmos w=1u l=1u
M11455 n4509 net3427 VSS VSS nmos w=1u l=1u
M11456 net3427 n4430 net3428 VSS nmos w=1u l=1u
M11457 net3427 net3425 net3426 VSS nmos w=1u l=1u
M11458 net3428 net3426 VSS VSS nmos w=1u l=1u
M11459 net3427 net3425 net3429 VDD pmos w=2u l=1u
M11460 net3425 n4430 VDD VDD pmos w=2u l=1u
M11461 net3426 n4430 net3427 VDD pmos w=2u l=1u
M11462 net3426 n4431 VDD VDD pmos w=2u l=1u
M11463 n4509 net3427 VDD VDD pmos w=2u l=1u
M11464 net3429 net3426 VDD VDD pmos w=2u l=1u
M11465 n4430 n4504 VDD VDD pmos w=2u l=1u
M11466 n4430 n4504 VSS VSS nmos w=1u l=1u
M11467 n4508 n4516 net3430 VSS nmos w=1u l=1u
M11468 net3430 n4515 VSS VSS nmos w=1u l=1u
M11469 n4508 n4516 VDD VDD pmos w=2u l=1u
M11470 n4508 n4515 VDD VDD pmos w=2u l=1u
M11471 net3431 n4431 VSS VSS nmos w=1u l=1u
M11472 net3432 n4504 VSS VSS nmos w=1u l=1u
M11473 n4516 net3433 VSS VSS nmos w=1u l=1u
M11474 net3433 n4431 net3434 VSS nmos w=1u l=1u
M11475 net3433 net3431 net3432 VSS nmos w=1u l=1u
M11476 net3434 net3432 VSS VSS nmos w=1u l=1u
M11477 net3433 net3431 net3435 VDD pmos w=2u l=1u
M11478 net3431 n4431 VDD VDD pmos w=2u l=1u
M11479 net3432 n4431 net3433 VDD pmos w=2u l=1u
M11480 net3432 n4504 VDD VDD pmos w=2u l=1u
M11481 n4516 net3433 VDD VDD pmos w=2u l=1u
M11482 net3435 net3432 VDD VDD pmos w=2u l=1u
M11483 n4431 N392 net3436 VSS nmos w=1u l=1u
M11484 net3436 N18 VSS VSS nmos w=1u l=1u
M11485 n4431 N392 VDD VDD pmos w=2u l=1u
M11486 n4431 N18 VDD VDD pmos w=2u l=1u
M11487 n4504 n4429 net3437 VSS nmos w=1u l=1u
M11488 net3437 n4517 VSS VSS nmos w=1u l=1u
M11489 n4504 n4429 VDD VDD pmos w=2u l=1u
M11490 n4504 n4517 VDD VDD pmos w=2u l=1u
M11491 n4429 n4519 net3438 VSS nmos w=1u l=1u
M11492 net3438 n4518 VSS VSS nmos w=1u l=1u
M11493 n4429 n4519 VDD VDD pmos w=2u l=1u
M11494 n4429 n4518 VDD VDD pmos w=2u l=1u
M11495 n4519 n4521 net3439 VSS nmos w=1u l=1u
M11496 net3439 n4520 VSS VSS nmos w=1u l=1u
M11497 n4519 n4521 VDD VDD pmos w=2u l=1u
M11498 n4519 n4520 VDD VDD pmos w=2u l=1u
M11499 n4520 n4523 net3440 VSS nmos w=1u l=1u
M11500 net3440 n4522 VSS VSS nmos w=1u l=1u
M11501 n4520 n4523 VDD VDD pmos w=2u l=1u
M11502 n4520 n4522 VDD VDD pmos w=2u l=1u
M11503 net3441 n4439 VSS VSS nmos w=1u l=1u
M11504 net3442 n4440 VSS VSS nmos w=1u l=1u
M11505 n4518 net3443 VSS VSS nmos w=1u l=1u
M11506 net3443 n4439 net3444 VSS nmos w=1u l=1u
M11507 net3443 net3441 net3442 VSS nmos w=1u l=1u
M11508 net3444 net3442 VSS VSS nmos w=1u l=1u
M11509 net3443 net3441 net3445 VDD pmos w=2u l=1u
M11510 net3441 n4439 VDD VDD pmos w=2u l=1u
M11511 net3442 n4439 net3443 VDD pmos w=2u l=1u
M11512 net3442 n4440 VDD VDD pmos w=2u l=1u
M11513 n4518 net3443 VDD VDD pmos w=2u l=1u
M11514 net3445 net3442 VDD VDD pmos w=2u l=1u
M11515 n4439 n4500 VDD VDD pmos w=2u l=1u
M11516 n4439 n4500 VSS VSS nmos w=1u l=1u
M11517 n4517 n4525 net3446 VSS nmos w=1u l=1u
M11518 net3446 n4524 VSS VSS nmos w=1u l=1u
M11519 n4517 n4525 VDD VDD pmos w=2u l=1u
M11520 n4517 n4524 VDD VDD pmos w=2u l=1u
M11521 net3447 n4440 VSS VSS nmos w=1u l=1u
M11522 net3448 n4500 VSS VSS nmos w=1u l=1u
M11523 n4525 net3449 VSS VSS nmos w=1u l=1u
M11524 net3449 n4440 net3450 VSS nmos w=1u l=1u
M11525 net3449 net3447 net3448 VSS nmos w=1u l=1u
M11526 net3450 net3448 VSS VSS nmos w=1u l=1u
M11527 net3449 net3447 net3451 VDD pmos w=2u l=1u
M11528 net3447 n4440 VDD VDD pmos w=2u l=1u
M11529 net3448 n4440 net3449 VDD pmos w=2u l=1u
M11530 net3448 n4500 VDD VDD pmos w=2u l=1u
M11531 n4525 net3449 VDD VDD pmos w=2u l=1u
M11532 net3451 net3448 VDD VDD pmos w=2u l=1u
M11533 n4440 N375 net3452 VSS nmos w=1u l=1u
M11534 net3452 N35 VSS VSS nmos w=1u l=1u
M11535 n4440 N375 VDD VDD pmos w=2u l=1u
M11536 n4440 N35 VDD VDD pmos w=2u l=1u
M11537 n4500 n4438 net3453 VSS nmos w=1u l=1u
M11538 net3453 n4526 VSS VSS nmos w=1u l=1u
M11539 n4500 n4438 VDD VDD pmos w=2u l=1u
M11540 n4500 n4526 VDD VDD pmos w=2u l=1u
M11541 n4438 n4528 net3454 VSS nmos w=1u l=1u
M11542 net3454 n4527 VSS VSS nmos w=1u l=1u
M11543 n4438 n4528 VDD VDD pmos w=2u l=1u
M11544 n4438 n4527 VDD VDD pmos w=2u l=1u
M11545 n4528 n4530 net3455 VSS nmos w=1u l=1u
M11546 net3455 n4529 VSS VSS nmos w=1u l=1u
M11547 n4528 n4530 VDD VDD pmos w=2u l=1u
M11548 n4528 n4529 VDD VDD pmos w=2u l=1u
M11549 n4529 net3456 VSS VSS nmos w=1u l=1u
M11550 net3456 n4531 VSS VSS nmos w=1u l=1u
M11551 net3456 n4532 VSS VSS nmos w=1u l=1u
M11552 net3456 n4532 net3457 VDD pmos w=2u l=1u
M11553 n4529 net3456 VDD VDD pmos w=2u l=1u
M11554 net3457 n4531 VDD VDD pmos w=2u l=1u
M11555 net3458 n4449 VSS VSS nmos w=1u l=1u
M11556 net3459 n4450 VSS VSS nmos w=1u l=1u
M11557 n4527 net3460 VSS VSS nmos w=1u l=1u
M11558 net3460 n4449 net3461 VSS nmos w=1u l=1u
M11559 net3460 net3458 net3459 VSS nmos w=1u l=1u
M11560 net3461 net3459 VSS VSS nmos w=1u l=1u
M11561 net3460 net3458 net3462 VDD pmos w=2u l=1u
M11562 net3458 n4449 VDD VDD pmos w=2u l=1u
M11563 net3459 n4449 net3460 VDD pmos w=2u l=1u
M11564 net3459 n4450 VDD VDD pmos w=2u l=1u
M11565 n4527 net3460 VDD VDD pmos w=2u l=1u
M11566 net3462 net3459 VDD VDD pmos w=2u l=1u
M11567 n4450 n4533 VDD VDD pmos w=2u l=1u
M11568 n4450 n4533 VSS VSS nmos w=1u l=1u
M11569 n4526 n4535 net3463 VSS nmos w=1u l=1u
M11570 net3463 n4534 VSS VSS nmos w=1u l=1u
M11571 n4526 n4535 VDD VDD pmos w=2u l=1u
M11572 n4526 n4534 VDD VDD pmos w=2u l=1u
M11573 net3464 n4533 VSS VSS nmos w=1u l=1u
M11574 net3465 n4449 VSS VSS nmos w=1u l=1u
M11575 n4535 net3466 VSS VSS nmos w=1u l=1u
M11576 net3466 n4533 net3467 VSS nmos w=1u l=1u
M11577 net3466 net3464 net3465 VSS nmos w=1u l=1u
M11578 net3467 net3465 VSS VSS nmos w=1u l=1u
M11579 net3466 net3464 net3468 VDD pmos w=2u l=1u
M11580 net3464 n4533 VDD VDD pmos w=2u l=1u
M11581 net3465 n4533 net3466 VDD pmos w=2u l=1u
M11582 net3465 n4449 VDD VDD pmos w=2u l=1u
M11583 n4535 net3466 VDD VDD pmos w=2u l=1u
M11584 net3468 net3465 VDD VDD pmos w=2u l=1u
M11585 n4533 N358 net3469 VSS nmos w=1u l=1u
M11586 net3469 N52 VSS VSS nmos w=1u l=1u
M11587 n4533 N358 VDD VDD pmos w=2u l=1u
M11588 n4533 N52 VDD VDD pmos w=2u l=1u
M11589 n4449 n4448 net3470 VSS nmos w=1u l=1u
M11590 net3470 n4536 VSS VSS nmos w=1u l=1u
M11591 n4449 n4448 VDD VDD pmos w=2u l=1u
M11592 n4449 n4536 VDD VDD pmos w=2u l=1u
M11593 n4448 n4538 net3471 VSS nmos w=1u l=1u
M11594 net3471 n4537 VSS VSS nmos w=1u l=1u
M11595 n4448 n4538 VDD VDD pmos w=2u l=1u
M11596 n4448 n4537 VDD VDD pmos w=2u l=1u
M11597 n4538 n4540 net3472 VSS nmos w=1u l=1u
M11598 net3472 n4539 VSS VSS nmos w=1u l=1u
M11599 n4538 n4540 VDD VDD pmos w=2u l=1u
M11600 n4538 n4539 VDD VDD pmos w=2u l=1u
M11601 n4539 n4542 net3473 VSS nmos w=1u l=1u
M11602 net3473 n4541 VSS VSS nmos w=1u l=1u
M11603 n4539 n4542 VDD VDD pmos w=2u l=1u
M11604 n4539 n4541 VDD VDD pmos w=2u l=1u
M11605 net3474 n4459 VSS VSS nmos w=1u l=1u
M11606 net3475 n4460 VSS VSS nmos w=1u l=1u
M11607 n4537 net3476 VSS VSS nmos w=1u l=1u
M11608 net3476 n4459 net3477 VSS nmos w=1u l=1u
M11609 net3476 net3474 net3475 VSS nmos w=1u l=1u
M11610 net3477 net3475 VSS VSS nmos w=1u l=1u
M11611 net3476 net3474 net3478 VDD pmos w=2u l=1u
M11612 net3474 n4459 VDD VDD pmos w=2u l=1u
M11613 net3475 n4459 net3476 VDD pmos w=2u l=1u
M11614 net3475 n4460 VDD VDD pmos w=2u l=1u
M11615 n4537 net3476 VDD VDD pmos w=2u l=1u
M11616 net3478 net3475 VDD VDD pmos w=2u l=1u
M11617 n4459 n4543 VDD VDD pmos w=2u l=1u
M11618 n4459 n4543 VSS VSS nmos w=1u l=1u
M11619 n4536 n4545 net3479 VSS nmos w=1u l=1u
M11620 net3479 n4544 VSS VSS nmos w=1u l=1u
M11621 n4536 n4545 VDD VDD pmos w=2u l=1u
M11622 n4536 n4544 VDD VDD pmos w=2u l=1u
M11623 net3480 n4460 VSS VSS nmos w=1u l=1u
M11624 net3481 n4543 VSS VSS nmos w=1u l=1u
M11625 n4545 net3482 VSS VSS nmos w=1u l=1u
M11626 net3482 n4460 net3483 VSS nmos w=1u l=1u
M11627 net3482 net3480 net3481 VSS nmos w=1u l=1u
M11628 net3483 net3481 VSS VSS nmos w=1u l=1u
M11629 net3482 net3480 net3484 VDD pmos w=2u l=1u
M11630 net3480 n4460 VDD VDD pmos w=2u l=1u
M11631 net3481 n4460 net3482 VDD pmos w=2u l=1u
M11632 net3481 n4543 VDD VDD pmos w=2u l=1u
M11633 n4545 net3482 VDD VDD pmos w=2u l=1u
M11634 net3484 net3481 VDD VDD pmos w=2u l=1u
M11635 n4460 N341 net3485 VSS nmos w=1u l=1u
M11636 net3485 N69 VSS VSS nmos w=1u l=1u
M11637 n4460 N341 VDD VDD pmos w=2u l=1u
M11638 n4460 N69 VDD VDD pmos w=2u l=1u
M11639 n4543 n4458 net3486 VSS nmos w=1u l=1u
M11640 net3486 n4546 VSS VSS nmos w=1u l=1u
M11641 n4543 n4458 VDD VDD pmos w=2u l=1u
M11642 n4543 n4546 VDD VDD pmos w=2u l=1u
M11643 n4458 n4548 net3487 VSS nmos w=1u l=1u
M11644 net3487 n4547 VSS VSS nmos w=1u l=1u
M11645 n4458 n4548 VDD VDD pmos w=2u l=1u
M11646 n4458 n4547 VDD VDD pmos w=2u l=1u
M11647 n4548 net3488 VSS VSS nmos w=1u l=1u
M11648 net3488 n4549 VSS VSS nmos w=1u l=1u
M11649 net3488 n4550 VSS VSS nmos w=1u l=1u
M11650 net3488 n4550 net3489 VDD pmos w=2u l=1u
M11651 n4548 net3488 VDD VDD pmos w=2u l=1u
M11652 net3489 n4549 VDD VDD pmos w=2u l=1u
M11653 n4547 net3490 VSS VSS nmos w=1u l=1u
M11654 net3491 n4551 VSS VSS nmos w=1u l=1u
M11655 net3490 n4492 net3491 VSS nmos w=1u l=1u
M11656 net3490 n4551 VDD VDD pmos w=2u l=1u
M11657 net3490 n4492 VDD VDD pmos w=2u l=1u
M11658 n4547 net3490 VDD VDD pmos w=2u l=1u
M11659 n4546 n4553 net3492 VSS nmos w=1u l=1u
M11660 net3492 n4552 VSS VSS nmos w=1u l=1u
M11661 n4546 n4553 VDD VDD pmos w=2u l=1u
M11662 n4546 n4552 VDD VDD pmos w=2u l=1u
M11663 n4553 n4492 net3493 VSS nmos w=1u l=1u
M11664 net3493 n4551 VSS VSS nmos w=1u l=1u
M11665 n4553 n4492 VDD VDD pmos w=2u l=1u
M11666 n4553 n4551 VDD VDD pmos w=2u l=1u
M11667 n4492 n4555 net3494 VSS nmos w=1u l=1u
M11668 net3494 n4554 VSS VSS nmos w=1u l=1u
M11669 n4492 n4555 VDD VDD pmos w=2u l=1u
M11670 n4492 n4554 VDD VDD pmos w=2u l=1u
M11671 n4555 N324 net3495 VSS nmos w=1u l=1u
M11672 net3495 N86 VSS VSS nmos w=1u l=1u
M11673 n4555 N324 VDD VDD pmos w=2u l=1u
M11674 n4555 N86 VDD VDD pmos w=2u l=1u
M11675 n4551 N86 net3496 VSS nmos w=1u l=1u
M11676 net3496 n4556 VSS VSS nmos w=1u l=1u
M11677 n4551 N86 VDD VDD pmos w=2u l=1u
M11678 n4551 n4556 VDD VDD pmos w=2u l=1u
M11679 n4556 n3257 VSS VSS nmos w=1u l=1u
M11680 n4556 n4554 VSS VSS nmos w=1u l=1u
M11681 n4556 n3257 net3497 VDD pmos w=2u l=1u
M11682 net3497 n4554 VDD VDD pmos w=2u l=1u
M11683 n4554 n4468 VSS VSS nmos w=1u l=1u
M11684 n4554 n4557 VSS VSS nmos w=1u l=1u
M11685 n4554 n4468 net3498 VDD pmos w=2u l=1u
M11686 net3498 n4557 VDD VDD pmos w=2u l=1u
M11687 n4468 n4559 VSS VSS nmos w=1u l=1u
M11688 n4468 n4558 VSS VSS nmos w=1u l=1u
M11689 n4468 n4559 net3499 VDD pmos w=2u l=1u
M11690 net3499 n4558 VDD VDD pmos w=2u l=1u
M11691 n4557 net3500 VSS VSS nmos w=1u l=1u
M11692 net3501 n4558 VSS VSS nmos w=1u l=1u
M11693 net3500 n4559 net3501 VSS nmos w=1u l=1u
M11694 net3500 n4558 VDD VDD pmos w=2u l=1u
M11695 net3500 n4559 VDD VDD pmos w=2u l=1u
M11696 n4557 net3500 VDD VDD pmos w=2u l=1u
M11697 n4558 n4560 net3502 VSS nmos w=1u l=1u
M11698 net3502 n4490 VSS VSS nmos w=1u l=1u
M11699 n4558 n4560 VDD VDD pmos w=2u l=1u
M11700 n4558 n4490 VDD VDD pmos w=2u l=1u
M11701 n4560 N103 net3503 VSS nmos w=1u l=1u
M11702 net3503 n4561 VSS VSS nmos w=1u l=1u
M11703 n4560 N103 VDD VDD pmos w=2u l=1u
M11704 n4560 n4561 VDD VDD pmos w=2u l=1u
M11705 n4561 n3411 VSS VSS nmos w=1u l=1u
M11706 n4561 n4562 VSS VSS nmos w=1u l=1u
M11707 n4561 n3411 net3504 VDD pmos w=2u l=1u
M11708 net3504 n4562 VDD VDD pmos w=2u l=1u
M11709 n4490 n4563 net3505 VSS nmos w=1u l=1u
M11710 net3505 n4562 VSS VSS nmos w=1u l=1u
M11711 n4490 n4563 VDD VDD pmos w=2u l=1u
M11712 n4490 n4562 VDD VDD pmos w=2u l=1u
M11713 n4563 N307 net3506 VSS nmos w=1u l=1u
M11714 net3506 N103 VSS VSS nmos w=1u l=1u
M11715 n4563 N307 VDD VDD pmos w=2u l=1u
M11716 n4563 N103 VDD VDD pmos w=2u l=1u
M11717 n4562 net3507 VSS VSS nmos w=1u l=1u
M11718 net3508 n4564 VSS VSS nmos w=1u l=1u
M11719 net3507 n4491 net3508 VSS nmos w=1u l=1u
M11720 net3507 n4564 VDD VDD pmos w=2u l=1u
M11721 net3507 n4491 VDD VDD pmos w=2u l=1u
M11722 n4562 net3507 VDD VDD pmos w=2u l=1u
M11723 n4564 net3509 VSS VSS nmos w=1u l=1u
M11724 net3509 n4565 VSS VSS nmos w=1u l=1u
M11725 net3509 n4483 VSS VSS nmos w=1u l=1u
M11726 net3509 n4483 net3510 VDD pmos w=2u l=1u
M11727 n4564 net3509 VDD VDD pmos w=2u l=1u
M11728 net3510 n4565 VDD VDD pmos w=2u l=1u
M11729 n4483 n4484 VDD VDD pmos w=2u l=1u
M11730 n4483 n4484 VSS VSS nmos w=1u l=1u
M11731 n4491 n4566 net3511 VSS nmos w=1u l=1u
M11732 net3511 n4565 VSS VSS nmos w=1u l=1u
M11733 n4491 n4566 VDD VDD pmos w=2u l=1u
M11734 n4491 n4565 VDD VDD pmos w=2u l=1u
M11735 n4566 n4484 net3512 VSS nmos w=1u l=1u
M11736 net3512 n4567 VSS VSS nmos w=1u l=1u
M11737 n4566 n4484 VDD VDD pmos w=2u l=1u
M11738 n4566 n4567 VDD VDD pmos w=2u l=1u
M11739 n4484 N137 net3513 VSS nmos w=1u l=1u
M11740 net3513 n4568 VSS VSS nmos w=1u l=1u
M11741 n4484 N137 VDD VDD pmos w=2u l=1u
M11742 n4484 n4568 VDD VDD pmos w=2u l=1u
M11743 n4568 net3514 VSS VSS nmos w=1u l=1u
M11744 net3515 N120 VSS VSS nmos w=1u l=1u
M11745 net3514 n3741 net3515 VSS nmos w=1u l=1u
M11746 net3514 N120 VDD VDD pmos w=2u l=1u
M11747 net3514 n3741 VDD VDD pmos w=2u l=1u
M11748 n4568 net3514 VDD VDD pmos w=2u l=1u
M11749 n4567 n4570 net3516 VSS nmos w=1u l=1u
M11750 net3516 n4569 VSS VSS nmos w=1u l=1u
M11751 n4567 n4570 VDD VDD pmos w=2u l=1u
M11752 n4567 n4569 VDD VDD pmos w=2u l=1u
M11753 n4570 N273 net3517 VSS nmos w=1u l=1u
M11754 net3517 N137 VSS VSS nmos w=1u l=1u
M11755 n4570 N273 VDD VDD pmos w=2u l=1u
M11756 n4570 N137 VDD VDD pmos w=2u l=1u
M11757 n4569 N290 net3518 VSS nmos w=1u l=1u
M11758 net3518 N120 VSS VSS nmos w=1u l=1u
M11759 n4569 N290 VDD VDD pmos w=2u l=1u
M11760 n4569 N120 VDD VDD pmos w=2u l=1u
M11761 n4559 net3519 VSS VSS nmos w=1u l=1u
M11762 net3520 n4572 VSS VSS nmos w=1u l=1u
M11763 net3519 n4571 net3520 VSS nmos w=1u l=1u
M11764 net3519 n4572 VDD VDD pmos w=2u l=1u
M11765 net3519 n4571 VDD VDD pmos w=2u l=1u
M11766 n4559 net3519 VDD VDD pmos w=2u l=1u
M11767 n4552 n4549 VSS VSS nmos w=1u l=1u
M11768 n4552 n4550 VSS VSS nmos w=1u l=1u
M11769 n4552 n4549 net3521 VDD pmos w=2u l=1u
M11770 net3521 n4550 VDD VDD pmos w=2u l=1u
M11771 n4549 n4573 VDD VDD pmos w=2u l=1u
M11772 n4549 n4573 VSS VSS nmos w=1u l=1u
M11773 n4544 n4575 VSS VSS nmos w=1u l=1u
M11774 n4544 n4574 VSS VSS nmos w=1u l=1u
M11775 n4544 n4575 net3522 VDD pmos w=2u l=1u
M11776 net3522 n4574 VDD VDD pmos w=2u l=1u
M11777 n4575 net3523 VSS VSS nmos w=1u l=1u
M11778 net3524 n4541 VSS VSS nmos w=1u l=1u
M11779 net3523 n4542 net3524 VSS nmos w=1u l=1u
M11780 net3523 n4541 VDD VDD pmos w=2u l=1u
M11781 net3523 n4542 VDD VDD pmos w=2u l=1u
M11782 n4575 net3523 VDD VDD pmos w=2u l=1u
M11783 n4574 n4540 VDD VDD pmos w=2u l=1u
M11784 n4574 n4540 VSS VSS nmos w=1u l=1u
M11785 n4534 n4577 VSS VSS nmos w=1u l=1u
M11786 n4534 n4576 VSS VSS nmos w=1u l=1u
M11787 n4534 n4577 net3525 VDD pmos w=2u l=1u
M11788 net3525 n4576 VDD VDD pmos w=2u l=1u
M11789 n4577 n4531 VSS VSS nmos w=1u l=1u
M11790 n4577 n4532 VSS VSS nmos w=1u l=1u
M11791 n4577 n4531 net3526 VDD pmos w=2u l=1u
M11792 net3526 n4532 VDD VDD pmos w=2u l=1u
M11793 n4576 n4530 VDD VDD pmos w=2u l=1u
M11794 n4576 n4530 VSS VSS nmos w=1u l=1u
M11795 n4524 n4579 VSS VSS nmos w=1u l=1u
M11796 n4524 n4578 VSS VSS nmos w=1u l=1u
M11797 n4524 n4579 net3527 VDD pmos w=2u l=1u
M11798 net3527 n4578 VDD VDD pmos w=2u l=1u
M11799 n4579 n4581 VSS VSS nmos w=1u l=1u
M11800 n4579 n4580 VSS VSS nmos w=1u l=1u
M11801 n4579 n4581 net3528 VDD pmos w=2u l=1u
M11802 net3528 n4580 VDD VDD pmos w=2u l=1u
M11803 n4580 n4523 VDD VDD pmos w=2u l=1u
M11804 n4580 n4523 VSS VSS nmos w=1u l=1u
M11805 n4578 n4521 VDD VDD pmos w=2u l=1u
M11806 n4578 n4521 VSS VSS nmos w=1u l=1u
M11807 n4515 n4583 VSS VSS nmos w=1u l=1u
M11808 n4515 n4582 VSS VSS nmos w=1u l=1u
M11809 n4515 n4583 net3529 VDD pmos w=2u l=1u
M11810 net3529 n4582 VDD VDD pmos w=2u l=1u
M11811 n4583 n4513 VSS VSS nmos w=1u l=1u
M11812 n4583 n4514 VSS VSS nmos w=1u l=1u
M11813 n4583 n4513 net3530 VDD pmos w=2u l=1u
M11814 net3530 n4514 VDD VDD pmos w=2u l=1u
M11815 n4582 n4512 VDD VDD pmos w=2u l=1u
M11816 n4582 n4512 VSS VSS nmos w=1u l=1u
M11817 net3531 n4514 VSS VSS nmos w=1u l=1u
M11818 net3532 n4584 VSS VSS nmos w=1u l=1u
M11819 N3552 net3533 VSS VSS nmos w=1u l=1u
M11820 net3533 n4514 net3534 VSS nmos w=1u l=1u
M11821 net3533 net3531 net3532 VSS nmos w=1u l=1u
M11822 net3534 net3532 VSS VSS nmos w=1u l=1u
M11823 net3533 net3531 net3535 VDD pmos w=2u l=1u
M11824 net3531 n4514 VDD VDD pmos w=2u l=1u
M11825 net3532 n4514 net3533 VDD pmos w=2u l=1u
M11826 net3532 n4584 VDD VDD pmos w=2u l=1u
M11827 N3552 net3533 VDD VDD pmos w=2u l=1u
M11828 net3535 net3532 VDD VDD pmos w=2u l=1u
M11829 n4514 n2721 VSS VSS nmos w=1u l=1u
M11830 n4514 n3929 VSS VSS nmos w=1u l=1u
M11831 n4514 n2721 net3536 VDD pmos w=2u l=1u
M11832 net3536 n3929 VDD VDD pmos w=2u l=1u
M11833 n2721 N392 VDD VDD pmos w=2u l=1u
M11834 n2721 N392 VSS VSS nmos w=1u l=1u
M11835 n4584 n4513 VDD VDD pmos w=2u l=1u
M11836 n4584 n4513 VSS VSS nmos w=1u l=1u
M11837 n4513 n4512 net3537 VSS nmos w=1u l=1u
M11838 net3537 n4585 VSS VSS nmos w=1u l=1u
M11839 n4513 n4512 VDD VDD pmos w=2u l=1u
M11840 n4513 n4585 VDD VDD pmos w=2u l=1u
M11841 n4512 n4587 net3538 VSS nmos w=1u l=1u
M11842 net3538 n4586 VSS VSS nmos w=1u l=1u
M11843 n4512 n4587 VDD VDD pmos w=2u l=1u
M11844 n4512 n4586 VDD VDD pmos w=2u l=1u
M11845 n4587 n4589 net3539 VSS nmos w=1u l=1u
M11846 net3539 n4588 VSS VSS nmos w=1u l=1u
M11847 n4587 n4589 VDD VDD pmos w=2u l=1u
M11848 n4587 n4588 VDD VDD pmos w=2u l=1u
M11849 n4588 net3540 VSS VSS nmos w=1u l=1u
M11850 net3540 n4590 VSS VSS nmos w=1u l=1u
M11851 net3540 n4591 VSS VSS nmos w=1u l=1u
M11852 net3540 n4591 net3541 VDD pmos w=2u l=1u
M11853 n4588 net3540 VDD VDD pmos w=2u l=1u
M11854 net3541 n4590 VDD VDD pmos w=2u l=1u
M11855 net3542 n4522 VSS VSS nmos w=1u l=1u
M11856 net3543 n4523 VSS VSS nmos w=1u l=1u
M11857 n4586 net3544 VSS VSS nmos w=1u l=1u
M11858 net3544 n4522 net3545 VSS nmos w=1u l=1u
M11859 net3544 net3542 net3543 VSS nmos w=1u l=1u
M11860 net3545 net3543 VSS VSS nmos w=1u l=1u
M11861 net3544 net3542 net3546 VDD pmos w=2u l=1u
M11862 net3542 n4522 VDD VDD pmos w=2u l=1u
M11863 net3543 n4522 net3544 VDD pmos w=2u l=1u
M11864 net3543 n4523 VDD VDD pmos w=2u l=1u
M11865 n4586 net3544 VDD VDD pmos w=2u l=1u
M11866 net3546 net3543 VDD VDD pmos w=2u l=1u
M11867 n4522 n4581 VDD VDD pmos w=2u l=1u
M11868 n4522 n4581 VSS VSS nmos w=1u l=1u
M11869 n4585 n4593 net3547 VSS nmos w=1u l=1u
M11870 net3547 n4592 VSS VSS nmos w=1u l=1u
M11871 n4585 n4593 VDD VDD pmos w=2u l=1u
M11872 n4585 n4592 VDD VDD pmos w=2u l=1u
M11873 net3548 n4523 VSS VSS nmos w=1u l=1u
M11874 net3549 n4581 VSS VSS nmos w=1u l=1u
M11875 n4593 net3550 VSS VSS nmos w=1u l=1u
M11876 net3550 n4523 net3551 VSS nmos w=1u l=1u
M11877 net3550 net3548 net3549 VSS nmos w=1u l=1u
M11878 net3551 net3549 VSS VSS nmos w=1u l=1u
M11879 net3550 net3548 net3552 VDD pmos w=2u l=1u
M11880 net3548 n4523 VDD VDD pmos w=2u l=1u
M11881 net3549 n4523 net3550 VDD pmos w=2u l=1u
M11882 net3549 n4581 VDD VDD pmos w=2u l=1u
M11883 n4593 net3550 VDD VDD pmos w=2u l=1u
M11884 net3552 net3549 VDD VDD pmos w=2u l=1u
M11885 n4523 N375 net3553 VSS nmos w=1u l=1u
M11886 net3553 N18 VSS VSS nmos w=1u l=1u
M11887 n4523 N375 VDD VDD pmos w=2u l=1u
M11888 n4523 N18 VDD VDD pmos w=2u l=1u
M11889 n4581 n4521 net3554 VSS nmos w=1u l=1u
M11890 net3554 n4594 VSS VSS nmos w=1u l=1u
M11891 n4581 n4521 VDD VDD pmos w=2u l=1u
M11892 n4581 n4594 VDD VDD pmos w=2u l=1u
M11893 n4521 n4596 net3555 VSS nmos w=1u l=1u
M11894 net3555 n4595 VSS VSS nmos w=1u l=1u
M11895 n4521 n4596 VDD VDD pmos w=2u l=1u
M11896 n4521 n4595 VDD VDD pmos w=2u l=1u
M11897 n4596 n4598 net3556 VSS nmos w=1u l=1u
M11898 net3556 n4597 VSS VSS nmos w=1u l=1u
M11899 n4596 n4598 VDD VDD pmos w=2u l=1u
M11900 n4596 n4597 VDD VDD pmos w=2u l=1u
M11901 n4597 net3557 VSS VSS nmos w=1u l=1u
M11902 net3557 n4599 VSS VSS nmos w=1u l=1u
M11903 net3557 n4600 VSS VSS nmos w=1u l=1u
M11904 net3557 n4600 net3558 VDD pmos w=2u l=1u
M11905 n4597 net3557 VDD VDD pmos w=2u l=1u
M11906 net3558 n4599 VDD VDD pmos w=2u l=1u
M11907 net3559 n4531 VSS VSS nmos w=1u l=1u
M11908 net3560 n4532 VSS VSS nmos w=1u l=1u
M11909 n4595 net3561 VSS VSS nmos w=1u l=1u
M11910 net3561 n4531 net3562 VSS nmos w=1u l=1u
M11911 net3561 net3559 net3560 VSS nmos w=1u l=1u
M11912 net3562 net3560 VSS VSS nmos w=1u l=1u
M11913 net3561 net3559 net3563 VDD pmos w=2u l=1u
M11914 net3559 n4531 VDD VDD pmos w=2u l=1u
M11915 net3560 n4531 net3561 VDD pmos w=2u l=1u
M11916 net3560 n4532 VDD VDD pmos w=2u l=1u
M11917 n4595 net3561 VDD VDD pmos w=2u l=1u
M11918 net3563 net3560 VDD VDD pmos w=2u l=1u
M11919 n4594 n4602 net3564 VSS nmos w=1u l=1u
M11920 net3564 n4601 VSS VSS nmos w=1u l=1u
M11921 n4594 n4602 VDD VDD pmos w=2u l=1u
M11922 n4594 n4601 VDD VDD pmos w=2u l=1u
M11923 net3565 n4532 VSS VSS nmos w=1u l=1u
M11924 net3566 n4603 VSS VSS nmos w=1u l=1u
M11925 n4602 net3567 VSS VSS nmos w=1u l=1u
M11926 net3567 n4532 net3568 VSS nmos w=1u l=1u
M11927 net3567 net3565 net3566 VSS nmos w=1u l=1u
M11928 net3568 net3566 VSS VSS nmos w=1u l=1u
M11929 net3567 net3565 net3569 VDD pmos w=2u l=1u
M11930 net3565 n4532 VDD VDD pmos w=2u l=1u
M11931 net3566 n4532 net3567 VDD pmos w=2u l=1u
M11932 net3566 n4603 VDD VDD pmos w=2u l=1u
M11933 n4602 net3567 VDD VDD pmos w=2u l=1u
M11934 net3569 net3566 VDD VDD pmos w=2u l=1u
M11935 n4532 n2965 VSS VSS nmos w=1u l=1u
M11936 n4532 n3456 VSS VSS nmos w=1u l=1u
M11937 n4532 n2965 net3570 VDD pmos w=2u l=1u
M11938 net3570 n3456 VDD VDD pmos w=2u l=1u
M11939 n4603 n4531 VDD VDD pmos w=2u l=1u
M11940 n4603 n4531 VSS VSS nmos w=1u l=1u
M11941 n4531 n4530 net3571 VSS nmos w=1u l=1u
M11942 net3571 n4604 VSS VSS nmos w=1u l=1u
M11943 n4531 n4530 VDD VDD pmos w=2u l=1u
M11944 n4531 n4604 VDD VDD pmos w=2u l=1u
M11945 n4530 n4606 net3572 VSS nmos w=1u l=1u
M11946 net3572 n4605 VSS VSS nmos w=1u l=1u
M11947 n4530 n4606 VDD VDD pmos w=2u l=1u
M11948 n4530 n4605 VDD VDD pmos w=2u l=1u
M11949 n4606 n4608 net3573 VSS nmos w=1u l=1u
M11950 net3573 n4607 VSS VSS nmos w=1u l=1u
M11951 n4606 n4608 VDD VDD pmos w=2u l=1u
M11952 n4606 n4607 VDD VDD pmos w=2u l=1u
M11953 n4607 n4610 net3574 VSS nmos w=1u l=1u
M11954 net3574 n4609 VSS VSS nmos w=1u l=1u
M11955 n4607 n4610 VDD VDD pmos w=2u l=1u
M11956 n4607 n4609 VDD VDD pmos w=2u l=1u
M11957 net3575 n4541 VSS VSS nmos w=1u l=1u
M11958 net3576 n4542 VSS VSS nmos w=1u l=1u
M11959 n4605 net3577 VSS VSS nmos w=1u l=1u
M11960 net3577 n4541 net3578 VSS nmos w=1u l=1u
M11961 net3577 net3575 net3576 VSS nmos w=1u l=1u
M11962 net3578 net3576 VSS VSS nmos w=1u l=1u
M11963 net3577 net3575 net3579 VDD pmos w=2u l=1u
M11964 net3575 n4541 VDD VDD pmos w=2u l=1u
M11965 net3576 n4541 net3577 VDD pmos w=2u l=1u
M11966 net3576 n4542 VDD VDD pmos w=2u l=1u
M11967 n4605 net3577 VDD VDD pmos w=2u l=1u
M11968 net3579 net3576 VDD VDD pmos w=2u l=1u
M11969 n4541 n4611 VDD VDD pmos w=2u l=1u
M11970 n4541 n4611 VSS VSS nmos w=1u l=1u
M11971 n4604 n4613 net3580 VSS nmos w=1u l=1u
M11972 net3580 n4612 VSS VSS nmos w=1u l=1u
M11973 n4604 n4613 VDD VDD pmos w=2u l=1u
M11974 n4604 n4612 VDD VDD pmos w=2u l=1u
M11975 net3581 n4542 VSS VSS nmos w=1u l=1u
M11976 net3582 n4611 VSS VSS nmos w=1u l=1u
M11977 n4613 net3583 VSS VSS nmos w=1u l=1u
M11978 net3583 n4542 net3584 VSS nmos w=1u l=1u
M11979 net3583 net3581 net3582 VSS nmos w=1u l=1u
M11980 net3584 net3582 VSS VSS nmos w=1u l=1u
M11981 net3583 net3581 net3585 VDD pmos w=2u l=1u
M11982 net3581 n4542 VDD VDD pmos w=2u l=1u
M11983 net3582 n4542 net3583 VDD pmos w=2u l=1u
M11984 net3582 n4611 VDD VDD pmos w=2u l=1u
M11985 n4613 net3583 VDD VDD pmos w=2u l=1u
M11986 net3585 net3582 VDD VDD pmos w=2u l=1u
M11987 n4542 N341 net3586 VSS nmos w=1u l=1u
M11988 net3586 N52 VSS VSS nmos w=1u l=1u
M11989 n4542 N341 VDD VDD pmos w=2u l=1u
M11990 n4542 N52 VDD VDD pmos w=2u l=1u
M11991 n4611 n4540 net3587 VSS nmos w=1u l=1u
M11992 net3587 n4614 VSS VSS nmos w=1u l=1u
M11993 n4611 n4540 VDD VDD pmos w=2u l=1u
M11994 n4611 n4614 VDD VDD pmos w=2u l=1u
M11995 n4540 n4616 net3588 VSS nmos w=1u l=1u
M11996 net3588 n4615 VSS VSS nmos w=1u l=1u
M11997 n4540 n4616 VDD VDD pmos w=2u l=1u
M11998 n4540 n4615 VDD VDD pmos w=2u l=1u
M11999 n4616 net3589 VSS VSS nmos w=1u l=1u
M12000 net3589 n4617 VSS VSS nmos w=1u l=1u
M12001 net3589 n4618 VSS VSS nmos w=1u l=1u
M12002 net3589 n4618 net3590 VDD pmos w=2u l=1u
M12003 n4616 net3589 VDD VDD pmos w=2u l=1u
M12004 net3590 n4617 VDD VDD pmos w=2u l=1u
M12005 n4615 net3591 VSS VSS nmos w=1u l=1u
M12006 net3592 n4619 VSS VSS nmos w=1u l=1u
M12007 net3591 n4573 net3592 VSS nmos w=1u l=1u
M12008 net3591 n4619 VDD VDD pmos w=2u l=1u
M12009 net3591 n4573 VDD VDD pmos w=2u l=1u
M12010 n4615 net3591 VDD VDD pmos w=2u l=1u
M12011 n4614 n4621 net3593 VSS nmos w=1u l=1u
M12012 net3593 n4620 VSS VSS nmos w=1u l=1u
M12013 n4614 n4621 VDD VDD pmos w=2u l=1u
M12014 n4614 n4620 VDD VDD pmos w=2u l=1u
M12015 n4621 n4573 net3594 VSS nmos w=1u l=1u
M12016 net3594 n4619 VSS VSS nmos w=1u l=1u
M12017 n4621 n4573 VDD VDD pmos w=2u l=1u
M12018 n4621 n4619 VDD VDD pmos w=2u l=1u
M12019 n4573 n4623 net3595 VSS nmos w=1u l=1u
M12020 net3595 n4622 VSS VSS nmos w=1u l=1u
M12021 n4573 n4623 VDD VDD pmos w=2u l=1u
M12022 n4573 n4622 VDD VDD pmos w=2u l=1u
M12023 n4623 N324 net3596 VSS nmos w=1u l=1u
M12024 net3596 N69 VSS VSS nmos w=1u l=1u
M12025 n4623 N324 VDD VDD pmos w=2u l=1u
M12026 n4623 N69 VDD VDD pmos w=2u l=1u
M12027 n4619 N69 net3597 VSS nmos w=1u l=1u
M12028 net3597 n4624 VSS VSS nmos w=1u l=1u
M12029 n4619 N69 VDD VDD pmos w=2u l=1u
M12030 n4619 n4624 VDD VDD pmos w=2u l=1u
M12031 n4624 n3257 VSS VSS nmos w=1u l=1u
M12032 n4624 n4622 VSS VSS nmos w=1u l=1u
M12033 n4624 n3257 net3598 VDD pmos w=2u l=1u
M12034 net3598 n4622 VDD VDD pmos w=2u l=1u
M12035 n4622 n4550 VSS VSS nmos w=1u l=1u
M12036 n4622 n4625 VSS VSS nmos w=1u l=1u
M12037 n4622 n4550 net3599 VDD pmos w=2u l=1u
M12038 net3599 n4625 VDD VDD pmos w=2u l=1u
M12039 n4550 n4627 VSS VSS nmos w=1u l=1u
M12040 n4550 n4626 VSS VSS nmos w=1u l=1u
M12041 n4550 n4627 net3600 VDD pmos w=2u l=1u
M12042 net3600 n4626 VDD VDD pmos w=2u l=1u
M12043 n4625 net3601 VSS VSS nmos w=1u l=1u
M12044 net3602 n4626 VSS VSS nmos w=1u l=1u
M12045 net3601 n4627 net3602 VSS nmos w=1u l=1u
M12046 net3601 n4626 VDD VDD pmos w=2u l=1u
M12047 net3601 n4627 VDD VDD pmos w=2u l=1u
M12048 n4625 net3601 VDD VDD pmos w=2u l=1u
M12049 n4626 n4628 net3603 VSS nmos w=1u l=1u
M12050 net3603 n4571 VSS VSS nmos w=1u l=1u
M12051 n4626 n4628 VDD VDD pmos w=2u l=1u
M12052 n4626 n4571 VDD VDD pmos w=2u l=1u
M12053 n4628 N86 net3604 VSS nmos w=1u l=1u
M12054 net3604 n4629 VSS VSS nmos w=1u l=1u
M12055 n4628 N86 VDD VDD pmos w=2u l=1u
M12056 n4628 n4629 VDD VDD pmos w=2u l=1u
M12057 n4629 n3411 VSS VSS nmos w=1u l=1u
M12058 n4629 n4630 VSS VSS nmos w=1u l=1u
M12059 n4629 n3411 net3605 VDD pmos w=2u l=1u
M12060 net3605 n4630 VDD VDD pmos w=2u l=1u
M12061 n4571 n4631 net3606 VSS nmos w=1u l=1u
M12062 net3606 n4630 VSS VSS nmos w=1u l=1u
M12063 n4571 n4631 VDD VDD pmos w=2u l=1u
M12064 n4571 n4630 VDD VDD pmos w=2u l=1u
M12065 n4631 N307 net3607 VSS nmos w=1u l=1u
M12066 net3607 N86 VSS VSS nmos w=1u l=1u
M12067 n4631 N307 VDD VDD pmos w=2u l=1u
M12068 n4631 N86 VDD VDD pmos w=2u l=1u
M12069 n4630 net3608 VSS VSS nmos w=1u l=1u
M12070 net3609 n4632 VSS VSS nmos w=1u l=1u
M12071 net3608 n4572 net3609 VSS nmos w=1u l=1u
M12072 net3608 n4632 VDD VDD pmos w=2u l=1u
M12073 net3608 n4572 VDD VDD pmos w=2u l=1u
M12074 n4630 net3608 VDD VDD pmos w=2u l=1u
M12075 n4632 n4565 net3610 VSS nmos w=1u l=1u
M12076 net3610 n4633 VSS VSS nmos w=1u l=1u
M12077 n4632 n4565 VDD VDD pmos w=2u l=1u
M12078 n4632 n4633 VDD VDD pmos w=2u l=1u
M12079 n4572 n4635 net3611 VSS nmos w=1u l=1u
M12080 net3611 n4634 VSS VSS nmos w=1u l=1u
M12081 n4572 n4635 VDD VDD pmos w=2u l=1u
M12082 n4572 n4634 VDD VDD pmos w=2u l=1u
M12083 n4635 n4565 net3612 VSS nmos w=1u l=1u
M12084 net3612 n4636 VSS VSS nmos w=1u l=1u
M12085 n4635 n4565 VDD VDD pmos w=2u l=1u
M12086 n4635 n4636 VDD VDD pmos w=2u l=1u
M12087 n4565 N120 net3613 VSS nmos w=1u l=1u
M12088 net3613 n4637 VSS VSS nmos w=1u l=1u
M12089 n4565 N120 VDD VDD pmos w=2u l=1u
M12090 n4565 n4637 VDD VDD pmos w=2u l=1u
M12091 n4637 net3614 VSS VSS nmos w=1u l=1u
M12092 net3615 N103 VSS VSS nmos w=1u l=1u
M12093 net3614 n3741 net3615 VSS nmos w=1u l=1u
M12094 net3614 N103 VDD VDD pmos w=2u l=1u
M12095 net3614 n3741 VDD VDD pmos w=2u l=1u
M12096 n4637 net3614 VDD VDD pmos w=2u l=1u
M12097 n4636 n4639 net3616 VSS nmos w=1u l=1u
M12098 net3616 n4638 VSS VSS nmos w=1u l=1u
M12099 n4636 n4639 VDD VDD pmos w=2u l=1u
M12100 n4636 n4638 VDD VDD pmos w=2u l=1u
M12101 n4639 N273 net3617 VSS nmos w=1u l=1u
M12102 net3617 N120 VSS VSS nmos w=1u l=1u
M12103 n4639 N273 VDD VDD pmos w=2u l=1u
M12104 n4639 N120 VDD VDD pmos w=2u l=1u
M12105 n4638 N290 net3618 VSS nmos w=1u l=1u
M12106 net3618 N103 VSS VSS nmos w=1u l=1u
M12107 n4638 N290 VDD VDD pmos w=2u l=1u
M12108 n4638 N103 VDD VDD pmos w=2u l=1u
M12109 n4627 net3619 VSS VSS nmos w=1u l=1u
M12110 net3620 n4641 VSS VSS nmos w=1u l=1u
M12111 net3619 n4640 net3620 VSS nmos w=1u l=1u
M12112 net3619 n4641 VDD VDD pmos w=2u l=1u
M12113 net3619 n4640 VDD VDD pmos w=2u l=1u
M12114 n4627 net3619 VDD VDD pmos w=2u l=1u
M12115 n4620 n4617 VSS VSS nmos w=1u l=1u
M12116 n4620 n4618 VSS VSS nmos w=1u l=1u
M12117 n4620 n4617 net3621 VDD pmos w=2u l=1u
M12118 net3621 n4618 VDD VDD pmos w=2u l=1u
M12119 n4617 n4642 VDD VDD pmos w=2u l=1u
M12120 n4617 n4642 VSS VSS nmos w=1u l=1u
M12121 n4612 n4644 VSS VSS nmos w=1u l=1u
M12122 n4612 n4643 VSS VSS nmos w=1u l=1u
M12123 n4612 n4644 net3622 VDD pmos w=2u l=1u
M12124 net3622 n4643 VDD VDD pmos w=2u l=1u
M12125 n4644 n4646 VSS VSS nmos w=1u l=1u
M12126 n4644 n4645 VSS VSS nmos w=1u l=1u
M12127 n4644 n4646 net3623 VDD pmos w=2u l=1u
M12128 net3623 n4645 VDD VDD pmos w=2u l=1u
M12129 n4645 n4610 VDD VDD pmos w=2u l=1u
M12130 n4645 n4610 VSS VSS nmos w=1u l=1u
M12131 n4643 n4608 VDD VDD pmos w=2u l=1u
M12132 n4643 n4608 VSS VSS nmos w=1u l=1u
M12133 n4601 n4648 VSS VSS nmos w=1u l=1u
M12134 n4601 n4647 VSS VSS nmos w=1u l=1u
M12135 n4601 n4648 net3624 VDD pmos w=2u l=1u
M12136 net3624 n4647 VDD VDD pmos w=2u l=1u
M12137 n4648 n4599 VSS VSS nmos w=1u l=1u
M12138 n4648 n4600 VSS VSS nmos w=1u l=1u
M12139 n4648 n4599 net3625 VDD pmos w=2u l=1u
M12140 net3625 n4600 VDD VDD pmos w=2u l=1u
M12141 n4647 n4598 VDD VDD pmos w=2u l=1u
M12142 n4647 n4598 VSS VSS nmos w=1u l=1u
M12143 n4592 n4650 VSS VSS nmos w=1u l=1u
M12144 n4592 n4649 VSS VSS nmos w=1u l=1u
M12145 n4592 n4650 net3626 VDD pmos w=2u l=1u
M12146 net3626 n4649 VDD VDD pmos w=2u l=1u
M12147 n4650 n4590 VSS VSS nmos w=1u l=1u
M12148 n4650 n4591 VSS VSS nmos w=1u l=1u
M12149 n4650 n4590 net3627 VDD pmos w=2u l=1u
M12150 net3627 n4591 VDD VDD pmos w=2u l=1u
M12151 n4649 n4589 VDD VDD pmos w=2u l=1u
M12152 n4649 n4589 VSS VSS nmos w=1u l=1u
M12153 net3628 n4591 VSS VSS nmos w=1u l=1u
M12154 net3629 n4651 VSS VSS nmos w=1u l=1u
M12155 N3211 net3630 VSS VSS nmos w=1u l=1u
M12156 net3630 n4591 net3631 VSS nmos w=1u l=1u
M12157 net3630 net3628 net3629 VSS nmos w=1u l=1u
M12158 net3631 net3629 VSS VSS nmos w=1u l=1u
M12159 net3630 net3628 net3632 VDD pmos w=2u l=1u
M12160 net3628 n4591 VDD VDD pmos w=2u l=1u
M12161 net3629 n4591 net3630 VDD pmos w=2u l=1u
M12162 net3629 n4651 VDD VDD pmos w=2u l=1u
M12163 N3211 net3630 VDD VDD pmos w=2u l=1u
M12164 net3632 net3629 VDD VDD pmos w=2u l=1u
M12165 n4591 n2837 VSS VSS nmos w=1u l=1u
M12166 n4591 n3929 VSS VSS nmos w=1u l=1u
M12167 n4591 n2837 net3633 VDD pmos w=2u l=1u
M12168 net3633 n3929 VDD VDD pmos w=2u l=1u
M12169 n2837 N375 VDD VDD pmos w=2u l=1u
M12170 n2837 N375 VSS VSS nmos w=1u l=1u
M12171 n4651 n4590 VDD VDD pmos w=2u l=1u
M12172 n4651 n4590 VSS VSS nmos w=1u l=1u
M12173 n4590 n4589 net3634 VSS nmos w=1u l=1u
M12174 net3634 n4652 VSS VSS nmos w=1u l=1u
M12175 n4590 n4589 VDD VDD pmos w=2u l=1u
M12176 n4590 n4652 VDD VDD pmos w=2u l=1u
M12177 n4589 n4654 net3635 VSS nmos w=1u l=1u
M12178 net3635 n4653 VSS VSS nmos w=1u l=1u
M12179 n4589 n4654 VDD VDD pmos w=2u l=1u
M12180 n4589 n4653 VDD VDD pmos w=2u l=1u
M12181 n4654 n4656 net3636 VSS nmos w=1u l=1u
M12182 net3636 n4655 VSS VSS nmos w=1u l=1u
M12183 n4654 n4656 VDD VDD pmos w=2u l=1u
M12184 n4654 n4655 VDD VDD pmos w=2u l=1u
M12185 n4655 net3637 VSS VSS nmos w=1u l=1u
M12186 net3637 n4657 VSS VSS nmos w=1u l=1u
M12187 net3637 n4658 VSS VSS nmos w=1u l=1u
M12188 net3637 n4658 net3638 VDD pmos w=2u l=1u
M12189 n4655 net3637 VDD VDD pmos w=2u l=1u
M12190 net3638 n4657 VDD VDD pmos w=2u l=1u
M12191 net3639 n4599 VSS VSS nmos w=1u l=1u
M12192 net3640 n4600 VSS VSS nmos w=1u l=1u
M12193 n4653 net3641 VSS VSS nmos w=1u l=1u
M12194 net3641 n4599 net3642 VSS nmos w=1u l=1u
M12195 net3641 net3639 net3640 VSS nmos w=1u l=1u
M12196 net3642 net3640 VSS VSS nmos w=1u l=1u
M12197 net3641 net3639 net3643 VDD pmos w=2u l=1u
M12198 net3639 n4599 VDD VDD pmos w=2u l=1u
M12199 net3640 n4599 net3641 VDD pmos w=2u l=1u
M12200 net3640 n4600 VDD VDD pmos w=2u l=1u
M12201 n4653 net3641 VDD VDD pmos w=2u l=1u
M12202 net3643 net3640 VDD VDD pmos w=2u l=1u
M12203 n4652 n4660 net3644 VSS nmos w=1u l=1u
M12204 net3644 n4659 VSS VSS nmos w=1u l=1u
M12205 n4652 n4660 VDD VDD pmos w=2u l=1u
M12206 n4652 n4659 VDD VDD pmos w=2u l=1u
M12207 net3645 n4600 VSS VSS nmos w=1u l=1u
M12208 net3646 n4661 VSS VSS nmos w=1u l=1u
M12209 n4660 net3647 VSS VSS nmos w=1u l=1u
M12210 net3647 n4600 net3648 VSS nmos w=1u l=1u
M12211 net3647 net3645 net3646 VSS nmos w=1u l=1u
M12212 net3648 net3646 VSS VSS nmos w=1u l=1u
M12213 net3647 net3645 net3649 VDD pmos w=2u l=1u
M12214 net3645 n4600 VDD VDD pmos w=2u l=1u
M12215 net3646 n4600 net3647 VDD pmos w=2u l=1u
M12216 net3646 n4661 VDD VDD pmos w=2u l=1u
M12217 n4660 net3647 VDD VDD pmos w=2u l=1u
M12218 net3649 net3646 VDD VDD pmos w=2u l=1u
M12219 n4600 n2965 VSS VSS nmos w=1u l=1u
M12220 n4600 n3603 VSS VSS nmos w=1u l=1u
M12221 n4600 n2965 net3650 VDD pmos w=2u l=1u
M12222 net3650 n3603 VDD VDD pmos w=2u l=1u
M12223 n4661 n4599 VDD VDD pmos w=2u l=1u
M12224 n4661 n4599 VSS VSS nmos w=1u l=1u
M12225 n4599 n4598 net3651 VSS nmos w=1u l=1u
M12226 net3651 n4662 VSS VSS nmos w=1u l=1u
M12227 n4599 n4598 VDD VDD pmos w=2u l=1u
M12228 n4599 n4662 VDD VDD pmos w=2u l=1u
M12229 n4598 n4664 net3652 VSS nmos w=1u l=1u
M12230 net3652 n4663 VSS VSS nmos w=1u l=1u
M12231 n4598 n4664 VDD VDD pmos w=2u l=1u
M12232 n4598 n4663 VDD VDD pmos w=2u l=1u
M12233 n4664 n4666 net3653 VSS nmos w=1u l=1u
M12234 net3653 n4665 VSS VSS nmos w=1u l=1u
M12235 n4664 n4666 VDD VDD pmos w=2u l=1u
M12236 n4664 n4665 VDD VDD pmos w=2u l=1u
M12237 n4665 n4668 net3654 VSS nmos w=1u l=1u
M12238 net3654 n4667 VSS VSS nmos w=1u l=1u
M12239 n4665 n4668 VDD VDD pmos w=2u l=1u
M12240 n4665 n4667 VDD VDD pmos w=2u l=1u
M12241 net3655 n4609 VSS VSS nmos w=1u l=1u
M12242 net3656 n4610 VSS VSS nmos w=1u l=1u
M12243 n4663 net3657 VSS VSS nmos w=1u l=1u
M12244 net3657 n4609 net3658 VSS nmos w=1u l=1u
M12245 net3657 net3655 net3656 VSS nmos w=1u l=1u
M12246 net3658 net3656 VSS VSS nmos w=1u l=1u
M12247 net3657 net3655 net3659 VDD pmos w=2u l=1u
M12248 net3655 n4609 VDD VDD pmos w=2u l=1u
M12249 net3656 n4609 net3657 VDD pmos w=2u l=1u
M12250 net3656 n4610 VDD VDD pmos w=2u l=1u
M12251 n4663 net3657 VDD VDD pmos w=2u l=1u
M12252 net3659 net3656 VDD VDD pmos w=2u l=1u
M12253 n4609 n4646 VDD VDD pmos w=2u l=1u
M12254 n4609 n4646 VSS VSS nmos w=1u l=1u
M12255 n4662 n4670 net3660 VSS nmos w=1u l=1u
M12256 net3660 n4669 VSS VSS nmos w=1u l=1u
M12257 n4662 n4670 VDD VDD pmos w=2u l=1u
M12258 n4662 n4669 VDD VDD pmos w=2u l=1u
M12259 net3661 n4610 VSS VSS nmos w=1u l=1u
M12260 net3662 n4646 VSS VSS nmos w=1u l=1u
M12261 n4670 net3663 VSS VSS nmos w=1u l=1u
M12262 net3663 n4610 net3664 VSS nmos w=1u l=1u
M12263 net3663 net3661 net3662 VSS nmos w=1u l=1u
M12264 net3664 net3662 VSS VSS nmos w=1u l=1u
M12265 net3663 net3661 net3665 VDD pmos w=2u l=1u
M12266 net3661 n4610 VDD VDD pmos w=2u l=1u
M12267 net3662 n4610 net3663 VDD pmos w=2u l=1u
M12268 net3662 n4646 VDD VDD pmos w=2u l=1u
M12269 n4670 net3663 VDD VDD pmos w=2u l=1u
M12270 net3665 net3662 VDD VDD pmos w=2u l=1u
M12271 n4610 N341 net3666 VSS nmos w=1u l=1u
M12272 net3666 N35 VSS VSS nmos w=1u l=1u
M12273 n4610 N341 VDD VDD pmos w=2u l=1u
M12274 n4610 N35 VDD VDD pmos w=2u l=1u
M12275 n4646 n4608 net3667 VSS nmos w=1u l=1u
M12276 net3667 n4671 VSS VSS nmos w=1u l=1u
M12277 n4646 n4608 VDD VDD pmos w=2u l=1u
M12278 n4646 n4671 VDD VDD pmos w=2u l=1u
M12279 n4608 n4673 net3668 VSS nmos w=1u l=1u
M12280 net3668 n4672 VSS VSS nmos w=1u l=1u
M12281 n4608 n4673 VDD VDD pmos w=2u l=1u
M12282 n4608 n4672 VDD VDD pmos w=2u l=1u
M12283 n4673 net3669 VSS VSS nmos w=1u l=1u
M12284 net3669 n4674 VSS VSS nmos w=1u l=1u
M12285 net3669 n4675 VSS VSS nmos w=1u l=1u
M12286 net3669 n4675 net3670 VDD pmos w=2u l=1u
M12287 n4673 net3669 VDD VDD pmos w=2u l=1u
M12288 net3670 n4674 VDD VDD pmos w=2u l=1u
M12289 n4672 net3671 VSS VSS nmos w=1u l=1u
M12290 net3672 n4676 VSS VSS nmos w=1u l=1u
M12291 net3671 n4642 net3672 VSS nmos w=1u l=1u
M12292 net3671 n4676 VDD VDD pmos w=2u l=1u
M12293 net3671 n4642 VDD VDD pmos w=2u l=1u
M12294 n4672 net3671 VDD VDD pmos w=2u l=1u
M12295 n4671 n4678 net3673 VSS nmos w=1u l=1u
M12296 net3673 n4677 VSS VSS nmos w=1u l=1u
M12297 n4671 n4678 VDD VDD pmos w=2u l=1u
M12298 n4671 n4677 VDD VDD pmos w=2u l=1u
M12299 n4678 n4642 net3674 VSS nmos w=1u l=1u
M12300 net3674 n4676 VSS VSS nmos w=1u l=1u
M12301 n4678 n4642 VDD VDD pmos w=2u l=1u
M12302 n4678 n4676 VDD VDD pmos w=2u l=1u
M12303 n4642 n4680 net3675 VSS nmos w=1u l=1u
M12304 net3675 n4679 VSS VSS nmos w=1u l=1u
M12305 n4642 n4680 VDD VDD pmos w=2u l=1u
M12306 n4642 n4679 VDD VDD pmos w=2u l=1u
M12307 n4680 N324 net3676 VSS nmos w=1u l=1u
M12308 net3676 N52 VSS VSS nmos w=1u l=1u
M12309 n4680 N324 VDD VDD pmos w=2u l=1u
M12310 n4680 N52 VDD VDD pmos w=2u l=1u
M12311 n4676 N52 net3677 VSS nmos w=1u l=1u
M12312 net3677 n4681 VSS VSS nmos w=1u l=1u
M12313 n4676 N52 VDD VDD pmos w=2u l=1u
M12314 n4676 n4681 VDD VDD pmos w=2u l=1u
M12315 n4681 n3257 VSS VSS nmos w=1u l=1u
M12316 n4681 n4679 VSS VSS nmos w=1u l=1u
M12317 n4681 n3257 net3678 VDD pmos w=2u l=1u
M12318 net3678 n4679 VDD VDD pmos w=2u l=1u
M12319 n4679 n4618 VSS VSS nmos w=1u l=1u
M12320 n4679 n4682 VSS VSS nmos w=1u l=1u
M12321 n4679 n4618 net3679 VDD pmos w=2u l=1u
M12322 net3679 n4682 VDD VDD pmos w=2u l=1u
M12323 n4618 n4684 VSS VSS nmos w=1u l=1u
M12324 n4618 n4683 VSS VSS nmos w=1u l=1u
M12325 n4618 n4684 net3680 VDD pmos w=2u l=1u
M12326 net3680 n4683 VDD VDD pmos w=2u l=1u
M12327 n4682 net3681 VSS VSS nmos w=1u l=1u
M12328 net3682 n4683 VSS VSS nmos w=1u l=1u
M12329 net3681 n4684 net3682 VSS nmos w=1u l=1u
M12330 net3681 n4683 VDD VDD pmos w=2u l=1u
M12331 net3681 n4684 VDD VDD pmos w=2u l=1u
M12332 n4682 net3681 VDD VDD pmos w=2u l=1u
M12333 n4683 n4685 net3683 VSS nmos w=1u l=1u
M12334 net3683 n4640 VSS VSS nmos w=1u l=1u
M12335 n4683 n4685 VDD VDD pmos w=2u l=1u
M12336 n4683 n4640 VDD VDD pmos w=2u l=1u
M12337 n4685 N69 net3684 VSS nmos w=1u l=1u
M12338 net3684 n4686 VSS VSS nmos w=1u l=1u
M12339 n4685 N69 VDD VDD pmos w=2u l=1u
M12340 n4685 n4686 VDD VDD pmos w=2u l=1u
M12341 n4686 n3411 VSS VSS nmos w=1u l=1u
M12342 n4686 n4687 VSS VSS nmos w=1u l=1u
M12343 n4686 n3411 net3685 VDD pmos w=2u l=1u
M12344 net3685 n4687 VDD VDD pmos w=2u l=1u
M12345 n4640 n4688 net3686 VSS nmos w=1u l=1u
M12346 net3686 n4687 VSS VSS nmos w=1u l=1u
M12347 n4640 n4688 VDD VDD pmos w=2u l=1u
M12348 n4640 n4687 VDD VDD pmos w=2u l=1u
M12349 n4688 N307 net3687 VSS nmos w=1u l=1u
M12350 net3687 N69 VSS VSS nmos w=1u l=1u
M12351 n4688 N307 VDD VDD pmos w=2u l=1u
M12352 n4688 N69 VDD VDD pmos w=2u l=1u
M12353 n4687 net3688 VSS VSS nmos w=1u l=1u
M12354 net3689 n4689 VSS VSS nmos w=1u l=1u
M12355 net3688 n4641 net3689 VSS nmos w=1u l=1u
M12356 net3688 n4689 VDD VDD pmos w=2u l=1u
M12357 net3688 n4641 VDD VDD pmos w=2u l=1u
M12358 n4687 net3688 VDD VDD pmos w=2u l=1u
M12359 n4689 net3690 VSS VSS nmos w=1u l=1u
M12360 net3690 n4690 VSS VSS nmos w=1u l=1u
M12361 net3690 n4633 VSS VSS nmos w=1u l=1u
M12362 net3690 n4633 net3691 VDD pmos w=2u l=1u
M12363 n4689 net3690 VDD VDD pmos w=2u l=1u
M12364 net3691 n4690 VDD VDD pmos w=2u l=1u
M12365 n4633 n4634 VDD VDD pmos w=2u l=1u
M12366 n4633 n4634 VSS VSS nmos w=1u l=1u
M12367 n4641 n4691 net3692 VSS nmos w=1u l=1u
M12368 net3692 n4690 VSS VSS nmos w=1u l=1u
M12369 n4641 n4691 VDD VDD pmos w=2u l=1u
M12370 n4641 n4690 VDD VDD pmos w=2u l=1u
M12371 n4691 n4634 net3693 VSS nmos w=1u l=1u
M12372 net3693 n4692 VSS VSS nmos w=1u l=1u
M12373 n4691 n4634 VDD VDD pmos w=2u l=1u
M12374 n4691 n4692 VDD VDD pmos w=2u l=1u
M12375 n4634 N103 net3694 VSS nmos w=1u l=1u
M12376 net3694 n4693 VSS VSS nmos w=1u l=1u
M12377 n4634 N103 VDD VDD pmos w=2u l=1u
M12378 n4634 n4693 VDD VDD pmos w=2u l=1u
M12379 n4693 net3695 VSS VSS nmos w=1u l=1u
M12380 net3696 N86 VSS VSS nmos w=1u l=1u
M12381 net3695 n3741 net3696 VSS nmos w=1u l=1u
M12382 net3695 N86 VDD VDD pmos w=2u l=1u
M12383 net3695 n3741 VDD VDD pmos w=2u l=1u
M12384 n4693 net3695 VDD VDD pmos w=2u l=1u
M12385 n4692 n4695 net3697 VSS nmos w=1u l=1u
M12386 net3697 n4694 VSS VSS nmos w=1u l=1u
M12387 n4692 n4695 VDD VDD pmos w=2u l=1u
M12388 n4692 n4694 VDD VDD pmos w=2u l=1u
M12389 n4695 N273 net3698 VSS nmos w=1u l=1u
M12390 net3698 N103 VSS VSS nmos w=1u l=1u
M12391 n4695 N273 VDD VDD pmos w=2u l=1u
M12392 n4695 N103 VDD VDD pmos w=2u l=1u
M12393 n4694 N290 net3699 VSS nmos w=1u l=1u
M12394 net3699 N86 VSS VSS nmos w=1u l=1u
M12395 n4694 N290 VDD VDD pmos w=2u l=1u
M12396 n4694 N86 VDD VDD pmos w=2u l=1u
M12397 n4684 net3700 VSS VSS nmos w=1u l=1u
M12398 net3701 n4697 VSS VSS nmos w=1u l=1u
M12399 net3700 n4696 net3701 VSS nmos w=1u l=1u
M12400 net3700 n4697 VDD VDD pmos w=2u l=1u
M12401 net3700 n4696 VDD VDD pmos w=2u l=1u
M12402 n4684 net3700 VDD VDD pmos w=2u l=1u
M12403 n4677 n4674 VSS VSS nmos w=1u l=1u
M12404 n4677 n4675 VSS VSS nmos w=1u l=1u
M12405 n4677 n4674 net3702 VDD pmos w=2u l=1u
M12406 net3702 n4675 VDD VDD pmos w=2u l=1u
M12407 n4674 n4698 VDD VDD pmos w=2u l=1u
M12408 n4674 n4698 VSS VSS nmos w=1u l=1u
M12409 n4669 n4700 VSS VSS nmos w=1u l=1u
M12410 n4669 n4699 VSS VSS nmos w=1u l=1u
M12411 n4669 n4700 net3703 VDD pmos w=2u l=1u
M12412 net3703 n4699 VDD VDD pmos w=2u l=1u
M12413 n4700 n4702 VSS VSS nmos w=1u l=1u
M12414 n4700 n4701 VSS VSS nmos w=1u l=1u
M12415 n4700 n4702 net3704 VDD pmos w=2u l=1u
M12416 net3704 n4701 VDD VDD pmos w=2u l=1u
M12417 n4701 n4668 VDD VDD pmos w=2u l=1u
M12418 n4701 n4668 VSS VSS nmos w=1u l=1u
M12419 n4699 n4666 VDD VDD pmos w=2u l=1u
M12420 n4699 n4666 VSS VSS nmos w=1u l=1u
M12421 n4659 n4704 VSS VSS nmos w=1u l=1u
M12422 n4659 n4703 VSS VSS nmos w=1u l=1u
M12423 n4659 n4704 net3705 VDD pmos w=2u l=1u
M12424 net3705 n4703 VDD VDD pmos w=2u l=1u
M12425 n4704 n4657 VSS VSS nmos w=1u l=1u
M12426 n4704 n4658 VSS VSS nmos w=1u l=1u
M12427 n4704 n4657 net3706 VDD pmos w=2u l=1u
M12428 net3706 n4658 VDD VDD pmos w=2u l=1u
M12429 n4703 n4656 VDD VDD pmos w=2u l=1u
M12430 n4703 n4656 VSS VSS nmos w=1u l=1u
M12431 net3707 n4658 VSS VSS nmos w=1u l=1u
M12432 net3708 n4705 VSS VSS nmos w=1u l=1u
M12433 N2877 net3709 VSS VSS nmos w=1u l=1u
M12434 net3709 n4658 net3710 VSS nmos w=1u l=1u
M12435 net3709 net3707 net3708 VSS nmos w=1u l=1u
M12436 net3710 net3708 VSS VSS nmos w=1u l=1u
M12437 net3709 net3707 net3711 VDD pmos w=2u l=1u
M12438 net3707 n4658 VDD VDD pmos w=2u l=1u
M12439 net3708 n4658 net3709 VDD pmos w=2u l=1u
M12440 net3708 n4705 VDD VDD pmos w=2u l=1u
M12441 N2877 net3709 VDD VDD pmos w=2u l=1u
M12442 net3711 net3708 VDD VDD pmos w=2u l=1u
M12443 n4658 n2965 VSS VSS nmos w=1u l=1u
M12444 n4658 n3929 VSS VSS nmos w=1u l=1u
M12445 n4658 n2965 net3712 VDD pmos w=2u l=1u
M12446 net3712 n3929 VDD VDD pmos w=2u l=1u
M12447 n2965 N358 VDD VDD pmos w=2u l=1u
M12448 n2965 N358 VSS VSS nmos w=1u l=1u
M12449 n4705 n4657 VDD VDD pmos w=2u l=1u
M12450 n4705 n4657 VSS VSS nmos w=1u l=1u
M12451 n4657 n4656 net3713 VSS nmos w=1u l=1u
M12452 net3713 n4706 VSS VSS nmos w=1u l=1u
M12453 n4657 n4656 VDD VDD pmos w=2u l=1u
M12454 n4657 n4706 VDD VDD pmos w=2u l=1u
M12455 n4656 n4708 net3714 VSS nmos w=1u l=1u
M12456 net3714 n4707 VSS VSS nmos w=1u l=1u
M12457 n4656 n4708 VDD VDD pmos w=2u l=1u
M12458 n4656 n4707 VDD VDD pmos w=2u l=1u
M12459 n4708 n4710 net3715 VSS nmos w=1u l=1u
M12460 net3715 n4709 VSS VSS nmos w=1u l=1u
M12461 n4708 n4710 VDD VDD pmos w=2u l=1u
M12462 n4708 n4709 VDD VDD pmos w=2u l=1u
M12463 n4709 net3716 VSS VSS nmos w=1u l=1u
M12464 net3716 n4711 VSS VSS nmos w=1u l=1u
M12465 net3716 n4712 VSS VSS nmos w=1u l=1u
M12466 net3716 n4712 net3717 VDD pmos w=2u l=1u
M12467 n4709 net3716 VDD VDD pmos w=2u l=1u
M12468 net3717 n4711 VDD VDD pmos w=2u l=1u
M12469 net3718 n4667 VSS VSS nmos w=1u l=1u
M12470 net3719 n4668 VSS VSS nmos w=1u l=1u
M12471 n4707 net3720 VSS VSS nmos w=1u l=1u
M12472 net3720 n4667 net3721 VSS nmos w=1u l=1u
M12473 net3720 net3718 net3719 VSS nmos w=1u l=1u
M12474 net3721 net3719 VSS VSS nmos w=1u l=1u
M12475 net3720 net3718 net3722 VDD pmos w=2u l=1u
M12476 net3718 n4667 VDD VDD pmos w=2u l=1u
M12477 net3719 n4667 net3720 VDD pmos w=2u l=1u
M12478 net3719 n4668 VDD VDD pmos w=2u l=1u
M12479 n4707 net3720 VDD VDD pmos w=2u l=1u
M12480 net3722 net3719 VDD VDD pmos w=2u l=1u
M12481 n4667 n4702 VDD VDD pmos w=2u l=1u
M12482 n4667 n4702 VSS VSS nmos w=1u l=1u
M12483 n4706 n4714 net3723 VSS nmos w=1u l=1u
M12484 net3723 n4713 VSS VSS nmos w=1u l=1u
M12485 n4706 n4714 VDD VDD pmos w=2u l=1u
M12486 n4706 n4713 VDD VDD pmos w=2u l=1u
M12487 net3724 n4668 VSS VSS nmos w=1u l=1u
M12488 net3725 n4702 VSS VSS nmos w=1u l=1u
M12489 n4714 net3726 VSS VSS nmos w=1u l=1u
M12490 net3726 n4668 net3727 VSS nmos w=1u l=1u
M12491 net3726 net3724 net3725 VSS nmos w=1u l=1u
M12492 net3727 net3725 VSS VSS nmos w=1u l=1u
M12493 net3726 net3724 net3728 VDD pmos w=2u l=1u
M12494 net3724 n4668 VDD VDD pmos w=2u l=1u
M12495 net3725 n4668 net3726 VDD pmos w=2u l=1u
M12496 net3725 n4702 VDD VDD pmos w=2u l=1u
M12497 n4714 net3726 VDD VDD pmos w=2u l=1u
M12498 net3728 net3725 VDD VDD pmos w=2u l=1u
M12499 n4668 N341 net3729 VSS nmos w=1u l=1u
M12500 net3729 N18 VSS VSS nmos w=1u l=1u
M12501 n4668 N341 VDD VDD pmos w=2u l=1u
M12502 n4668 N18 VDD VDD pmos w=2u l=1u
M12503 n4702 n4666 net3730 VSS nmos w=1u l=1u
M12504 net3730 n4715 VSS VSS nmos w=1u l=1u
M12505 n4702 n4666 VDD VDD pmos w=2u l=1u
M12506 n4702 n4715 VDD VDD pmos w=2u l=1u
M12507 n4666 n4717 net3731 VSS nmos w=1u l=1u
M12508 net3731 n4716 VSS VSS nmos w=1u l=1u
M12509 n4666 n4717 VDD VDD pmos w=2u l=1u
M12510 n4666 n4716 VDD VDD pmos w=2u l=1u
M12511 n4717 net3732 VSS VSS nmos w=1u l=1u
M12512 net3732 n4718 VSS VSS nmos w=1u l=1u
M12513 net3732 n4719 VSS VSS nmos w=1u l=1u
M12514 net3732 n4719 net3733 VDD pmos w=2u l=1u
M12515 n4717 net3732 VDD VDD pmos w=2u l=1u
M12516 net3733 n4718 VDD VDD pmos w=2u l=1u
M12517 n4716 net3734 VSS VSS nmos w=1u l=1u
M12518 net3735 n4720 VSS VSS nmos w=1u l=1u
M12519 net3734 n4698 net3735 VSS nmos w=1u l=1u
M12520 net3734 n4720 VDD VDD pmos w=2u l=1u
M12521 net3734 n4698 VDD VDD pmos w=2u l=1u
M12522 n4716 net3734 VDD VDD pmos w=2u l=1u
M12523 n4715 n4722 net3736 VSS nmos w=1u l=1u
M12524 net3736 n4721 VSS VSS nmos w=1u l=1u
M12525 n4715 n4722 VDD VDD pmos w=2u l=1u
M12526 n4715 n4721 VDD VDD pmos w=2u l=1u
M12527 n4722 n4698 net3737 VSS nmos w=1u l=1u
M12528 net3737 n4720 VSS VSS nmos w=1u l=1u
M12529 n4722 n4698 VDD VDD pmos w=2u l=1u
M12530 n4722 n4720 VDD VDD pmos w=2u l=1u
M12531 n4698 n4724 net3738 VSS nmos w=1u l=1u
M12532 net3738 n4723 VSS VSS nmos w=1u l=1u
M12533 n4698 n4724 VDD VDD pmos w=2u l=1u
M12534 n4698 n4723 VDD VDD pmos w=2u l=1u
M12535 n4724 N324 net3739 VSS nmos w=1u l=1u
M12536 net3739 N35 VSS VSS nmos w=1u l=1u
M12537 n4724 N324 VDD VDD pmos w=2u l=1u
M12538 n4724 N35 VDD VDD pmos w=2u l=1u
M12539 n4720 N35 net3740 VSS nmos w=1u l=1u
M12540 net3740 n4725 VSS VSS nmos w=1u l=1u
M12541 n4720 N35 VDD VDD pmos w=2u l=1u
M12542 n4720 n4725 VDD VDD pmos w=2u l=1u
M12543 n4725 n3257 VSS VSS nmos w=1u l=1u
M12544 n4725 n4723 VSS VSS nmos w=1u l=1u
M12545 n4725 n3257 net3741 VDD pmos w=2u l=1u
M12546 net3741 n4723 VDD VDD pmos w=2u l=1u
M12547 n4723 n4675 VSS VSS nmos w=1u l=1u
M12548 n4723 n4726 VSS VSS nmos w=1u l=1u
M12549 n4723 n4675 net3742 VDD pmos w=2u l=1u
M12550 net3742 n4726 VDD VDD pmos w=2u l=1u
M12551 n4675 n4728 VSS VSS nmos w=1u l=1u
M12552 n4675 n4727 VSS VSS nmos w=1u l=1u
M12553 n4675 n4728 net3743 VDD pmos w=2u l=1u
M12554 net3743 n4727 VDD VDD pmos w=2u l=1u
M12555 n4726 net3744 VSS VSS nmos w=1u l=1u
M12556 net3745 n4727 VSS VSS nmos w=1u l=1u
M12557 net3744 n4728 net3745 VSS nmos w=1u l=1u
M12558 net3744 n4727 VDD VDD pmos w=2u l=1u
M12559 net3744 n4728 VDD VDD pmos w=2u l=1u
M12560 n4726 net3744 VDD VDD pmos w=2u l=1u
M12561 n4727 n4729 net3746 VSS nmos w=1u l=1u
M12562 net3746 n4696 VSS VSS nmos w=1u l=1u
M12563 n4727 n4729 VDD VDD pmos w=2u l=1u
M12564 n4727 n4696 VDD VDD pmos w=2u l=1u
M12565 n4729 N52 net3747 VSS nmos w=1u l=1u
M12566 net3747 n4730 VSS VSS nmos w=1u l=1u
M12567 n4729 N52 VDD VDD pmos w=2u l=1u
M12568 n4729 n4730 VDD VDD pmos w=2u l=1u
M12569 n4730 n3411 VSS VSS nmos w=1u l=1u
M12570 n4730 n4731 VSS VSS nmos w=1u l=1u
M12571 n4730 n3411 net3748 VDD pmos w=2u l=1u
M12572 net3748 n4731 VDD VDD pmos w=2u l=1u
M12573 n4696 n4732 net3749 VSS nmos w=1u l=1u
M12574 net3749 n4731 VSS VSS nmos w=1u l=1u
M12575 n4696 n4732 VDD VDD pmos w=2u l=1u
M12576 n4696 n4731 VDD VDD pmos w=2u l=1u
M12577 n4732 N307 net3750 VSS nmos w=1u l=1u
M12578 net3750 N52 VSS VSS nmos w=1u l=1u
M12579 n4732 N307 VDD VDD pmos w=2u l=1u
M12580 n4732 N52 VDD VDD pmos w=2u l=1u
M12581 n4731 net3751 VSS VSS nmos w=1u l=1u
M12582 net3752 n4733 VSS VSS nmos w=1u l=1u
M12583 net3751 n4697 net3752 VSS nmos w=1u l=1u
M12584 net3751 n4733 VDD VDD pmos w=2u l=1u
M12585 net3751 n4697 VDD VDD pmos w=2u l=1u
M12586 n4731 net3751 VDD VDD pmos w=2u l=1u
M12587 n4733 n4690 net3753 VSS nmos w=1u l=1u
M12588 net3753 n4734 VSS VSS nmos w=1u l=1u
M12589 n4733 n4690 VDD VDD pmos w=2u l=1u
M12590 n4733 n4734 VDD VDD pmos w=2u l=1u
M12591 n4697 n4736 net3754 VSS nmos w=1u l=1u
M12592 net3754 n4735 VSS VSS nmos w=1u l=1u
M12593 n4697 n4736 VDD VDD pmos w=2u l=1u
M12594 n4697 n4735 VDD VDD pmos w=2u l=1u
M12595 n4736 n4690 net3755 VSS nmos w=1u l=1u
M12596 net3755 n4737 VSS VSS nmos w=1u l=1u
M12597 n4736 n4690 VDD VDD pmos w=2u l=1u
M12598 n4736 n4737 VDD VDD pmos w=2u l=1u
M12599 n4690 N86 net3756 VSS nmos w=1u l=1u
M12600 net3756 n4738 VSS VSS nmos w=1u l=1u
M12601 n4690 N86 VDD VDD pmos w=2u l=1u
M12602 n4690 n4738 VDD VDD pmos w=2u l=1u
M12603 n4738 net3757 VSS VSS nmos w=1u l=1u
M12604 net3758 N69 VSS VSS nmos w=1u l=1u
M12605 net3757 n3741 net3758 VSS nmos w=1u l=1u
M12606 net3757 N69 VDD VDD pmos w=2u l=1u
M12607 net3757 n3741 VDD VDD pmos w=2u l=1u
M12608 n4738 net3757 VDD VDD pmos w=2u l=1u
M12609 n4737 n4740 net3759 VSS nmos w=1u l=1u
M12610 net3759 n4739 VSS VSS nmos w=1u l=1u
M12611 n4737 n4740 VDD VDD pmos w=2u l=1u
M12612 n4737 n4739 VDD VDD pmos w=2u l=1u
M12613 n4740 N273 net3760 VSS nmos w=1u l=1u
M12614 net3760 N86 VSS VSS nmos w=1u l=1u
M12615 n4740 N273 VDD VDD pmos w=2u l=1u
M12616 n4740 N86 VDD VDD pmos w=2u l=1u
M12617 n4739 N290 net3761 VSS nmos w=1u l=1u
M12618 net3761 N69 VSS VSS nmos w=1u l=1u
M12619 n4739 N290 VDD VDD pmos w=2u l=1u
M12620 n4739 N69 VDD VDD pmos w=2u l=1u
M12621 n4728 net3762 VSS VSS nmos w=1u l=1u
M12622 net3763 n4742 VSS VSS nmos w=1u l=1u
M12623 net3762 n4741 net3763 VSS nmos w=1u l=1u
M12624 net3762 n4742 VDD VDD pmos w=2u l=1u
M12625 net3762 n4741 VDD VDD pmos w=2u l=1u
M12626 n4728 net3762 VDD VDD pmos w=2u l=1u
M12627 n4721 n4718 VSS VSS nmos w=1u l=1u
M12628 n4721 n4719 VSS VSS nmos w=1u l=1u
M12629 n4721 n4718 net3764 VDD pmos w=2u l=1u
M12630 net3764 n4719 VDD VDD pmos w=2u l=1u
M12631 n4718 n4743 VDD VDD pmos w=2u l=1u
M12632 n4718 n4743 VSS VSS nmos w=1u l=1u
M12633 n4713 n4745 VSS VSS nmos w=1u l=1u
M12634 n4713 n4744 VSS VSS nmos w=1u l=1u
M12635 n4713 n4745 net3765 VDD pmos w=2u l=1u
M12636 net3765 n4744 VDD VDD pmos w=2u l=1u
M12637 n4745 n4711 VSS VSS nmos w=1u l=1u
M12638 n4745 n4712 VSS VSS nmos w=1u l=1u
M12639 n4745 n4711 net3766 VDD pmos w=2u l=1u
M12640 net3766 n4712 VDD VDD pmos w=2u l=1u
M12641 n4744 n4710 VDD VDD pmos w=2u l=1u
M12642 n4744 n4710 VSS VSS nmos w=1u l=1u
M12643 net3767 n4712 VSS VSS nmos w=1u l=1u
M12644 net3768 n4746 VSS VSS nmos w=1u l=1u
M12645 N2548 net3769 VSS VSS nmos w=1u l=1u
M12646 net3769 n4712 net3770 VSS nmos w=1u l=1u
M12647 net3769 net3767 net3768 VSS nmos w=1u l=1u
M12648 net3770 net3768 VSS VSS nmos w=1u l=1u
M12649 net3769 net3767 net3771 VDD pmos w=2u l=1u
M12650 net3767 n4712 VDD VDD pmos w=2u l=1u
M12651 net3768 n4712 net3769 VDD pmos w=2u l=1u
M12652 net3768 n4746 VDD VDD pmos w=2u l=1u
M12653 N2548 net3769 VDD VDD pmos w=2u l=1u
M12654 net3771 net3768 VDD VDD pmos w=2u l=1u
M12655 n4712 n3105 VSS VSS nmos w=1u l=1u
M12656 n4712 n3929 VSS VSS nmos w=1u l=1u
M12657 n4712 n3105 net3772 VDD pmos w=2u l=1u
M12658 net3772 n3929 VDD VDD pmos w=2u l=1u
M12659 n3105 N341 VDD VDD pmos w=2u l=1u
M12660 n3105 N341 VSS VSS nmos w=1u l=1u
M12661 n4746 n4711 VDD VDD pmos w=2u l=1u
M12662 n4746 n4711 VSS VSS nmos w=1u l=1u
M12663 n4711 n4710 net3773 VSS nmos w=1u l=1u
M12664 net3773 n4747 VSS VSS nmos w=1u l=1u
M12665 n4711 n4710 VDD VDD pmos w=2u l=1u
M12666 n4711 n4747 VDD VDD pmos w=2u l=1u
M12667 n4710 n4749 net3774 VSS nmos w=1u l=1u
M12668 net3774 n4748 VSS VSS nmos w=1u l=1u
M12669 n4710 n4749 VDD VDD pmos w=2u l=1u
M12670 n4710 n4748 VDD VDD pmos w=2u l=1u
M12671 n4749 n4751 net3775 VSS nmos w=1u l=1u
M12672 net3775 n4750 VSS VSS nmos w=1u l=1u
M12673 n4749 n4751 VDD VDD pmos w=2u l=1u
M12674 n4749 n4750 VDD VDD pmos w=2u l=1u
M12675 n4748 net3776 VSS VSS nmos w=1u l=1u
M12676 net3777 n4752 VSS VSS nmos w=1u l=1u
M12677 net3776 n4743 net3777 VSS nmos w=1u l=1u
M12678 net3776 n4752 VDD VDD pmos w=2u l=1u
M12679 net3776 n4743 VDD VDD pmos w=2u l=1u
M12680 n4748 net3776 VDD VDD pmos w=2u l=1u
M12681 n4747 n4754 net3778 VSS nmos w=1u l=1u
M12682 net3778 n4753 VSS VSS nmos w=1u l=1u
M12683 n4747 n4754 VDD VDD pmos w=2u l=1u
M12684 n4747 n4753 VDD VDD pmos w=2u l=1u
M12685 n4754 n4743 net3779 VSS nmos w=1u l=1u
M12686 net3779 n4752 VSS VSS nmos w=1u l=1u
M12687 n4754 n4743 VDD VDD pmos w=2u l=1u
M12688 n4754 n4752 VDD VDD pmos w=2u l=1u
M12689 n4743 n4756 net3780 VSS nmos w=1u l=1u
M12690 net3780 n4755 VSS VSS nmos w=1u l=1u
M12691 n4743 n4756 VDD VDD pmos w=2u l=1u
M12692 n4743 n4755 VDD VDD pmos w=2u l=1u
M12693 n4756 N324 net3781 VSS nmos w=1u l=1u
M12694 net3781 N18 VSS VSS nmos w=1u l=1u
M12695 n4756 N324 VDD VDD pmos w=2u l=1u
M12696 n4756 N18 VDD VDD pmos w=2u l=1u
M12697 n4752 N18 net3782 VSS nmos w=1u l=1u
M12698 net3782 n4757 VSS VSS nmos w=1u l=1u
M12699 n4752 N18 VDD VDD pmos w=2u l=1u
M12700 n4752 n4757 VDD VDD pmos w=2u l=1u
M12701 n4757 n3257 VSS VSS nmos w=1u l=1u
M12702 n4757 n4755 VSS VSS nmos w=1u l=1u
M12703 n4757 n3257 net3783 VDD pmos w=2u l=1u
M12704 net3783 n4755 VDD VDD pmos w=2u l=1u
M12705 n4755 n4719 VSS VSS nmos w=1u l=1u
M12706 n4755 n4758 VSS VSS nmos w=1u l=1u
M12707 n4755 n4719 net3784 VDD pmos w=2u l=1u
M12708 net3784 n4758 VDD VDD pmos w=2u l=1u
M12709 n4719 n4760 VSS VSS nmos w=1u l=1u
M12710 n4719 n4759 VSS VSS nmos w=1u l=1u
M12711 n4719 n4760 net3785 VDD pmos w=2u l=1u
M12712 net3785 n4759 VDD VDD pmos w=2u l=1u
M12713 n4758 net3786 VSS VSS nmos w=1u l=1u
M12714 net3787 n4759 VSS VSS nmos w=1u l=1u
M12715 net3786 n4760 net3787 VSS nmos w=1u l=1u
M12716 net3786 n4759 VDD VDD pmos w=2u l=1u
M12717 net3786 n4760 VDD VDD pmos w=2u l=1u
M12718 n4758 net3786 VDD VDD pmos w=2u l=1u
M12719 n4759 n4761 net3788 VSS nmos w=1u l=1u
M12720 net3788 n4741 VSS VSS nmos w=1u l=1u
M12721 n4759 n4761 VDD VDD pmos w=2u l=1u
M12722 n4759 n4741 VDD VDD pmos w=2u l=1u
M12723 n4761 N35 net3789 VSS nmos w=1u l=1u
M12724 net3789 n4762 VSS VSS nmos w=1u l=1u
M12725 n4761 N35 VDD VDD pmos w=2u l=1u
M12726 n4761 n4762 VDD VDD pmos w=2u l=1u
M12727 n4762 n3411 VSS VSS nmos w=1u l=1u
M12728 n4762 n4763 VSS VSS nmos w=1u l=1u
M12729 n4762 n3411 net3790 VDD pmos w=2u l=1u
M12730 net3790 n4763 VDD VDD pmos w=2u l=1u
M12731 n4741 n4764 net3791 VSS nmos w=1u l=1u
M12732 net3791 n4763 VSS VSS nmos w=1u l=1u
M12733 n4741 n4764 VDD VDD pmos w=2u l=1u
M12734 n4741 n4763 VDD VDD pmos w=2u l=1u
M12735 n4764 N307 net3792 VSS nmos w=1u l=1u
M12736 net3792 N35 VSS VSS nmos w=1u l=1u
M12737 n4764 N307 VDD VDD pmos w=2u l=1u
M12738 n4764 N35 VDD VDD pmos w=2u l=1u
M12739 n4763 net3793 VSS VSS nmos w=1u l=1u
M12740 net3794 n4765 VSS VSS nmos w=1u l=1u
M12741 net3793 n4742 net3794 VSS nmos w=1u l=1u
M12742 net3793 n4765 VDD VDD pmos w=2u l=1u
M12743 net3793 n4742 VDD VDD pmos w=2u l=1u
M12744 n4763 net3793 VDD VDD pmos w=2u l=1u
M12745 n4765 net3795 VSS VSS nmos w=1u l=1u
M12746 net3795 n4766 VSS VSS nmos w=1u l=1u
M12747 net3795 n4734 VSS VSS nmos w=1u l=1u
M12748 net3795 n4734 net3796 VDD pmos w=2u l=1u
M12749 n4765 net3795 VDD VDD pmos w=2u l=1u
M12750 net3796 n4766 VDD VDD pmos w=2u l=1u
M12751 n4734 n4735 VDD VDD pmos w=2u l=1u
M12752 n4734 n4735 VSS VSS nmos w=1u l=1u
M12753 n4742 n4767 net3797 VSS nmos w=1u l=1u
M12754 net3797 n4766 VSS VSS nmos w=1u l=1u
M12755 n4742 n4767 VDD VDD pmos w=2u l=1u
M12756 n4742 n4766 VDD VDD pmos w=2u l=1u
M12757 n4767 n4735 net3798 VSS nmos w=1u l=1u
M12758 net3798 n4768 VSS VSS nmos w=1u l=1u
M12759 n4767 n4735 VDD VDD pmos w=2u l=1u
M12760 n4767 n4768 VDD VDD pmos w=2u l=1u
M12761 n4735 N69 net3799 VSS nmos w=1u l=1u
M12762 net3799 n4769 VSS VSS nmos w=1u l=1u
M12763 n4735 N69 VDD VDD pmos w=2u l=1u
M12764 n4735 n4769 VDD VDD pmos w=2u l=1u
M12765 n4769 net3800 VSS VSS nmos w=1u l=1u
M12766 net3801 N52 VSS VSS nmos w=1u l=1u
M12767 net3800 n3741 net3801 VSS nmos w=1u l=1u
M12768 net3800 N52 VDD VDD pmos w=2u l=1u
M12769 net3800 n3741 VDD VDD pmos w=2u l=1u
M12770 n4769 net3800 VDD VDD pmos w=2u l=1u
M12771 n4768 n4771 net3802 VSS nmos w=1u l=1u
M12772 net3802 n4770 VSS VSS nmos w=1u l=1u
M12773 n4768 n4771 VDD VDD pmos w=2u l=1u
M12774 n4768 n4770 VDD VDD pmos w=2u l=1u
M12775 n4771 N273 net3803 VSS nmos w=1u l=1u
M12776 net3803 N69 VSS VSS nmos w=1u l=1u
M12777 n4771 N273 VDD VDD pmos w=2u l=1u
M12778 n4771 N69 VDD VDD pmos w=2u l=1u
M12779 n4770 N290 net3804 VSS nmos w=1u l=1u
M12780 net3804 N52 VSS VSS nmos w=1u l=1u
M12781 n4770 N290 VDD VDD pmos w=2u l=1u
M12782 n4770 N52 VDD VDD pmos w=2u l=1u
M12783 n4760 net3805 VSS VSS nmos w=1u l=1u
M12784 net3806 n4773 VSS VSS nmos w=1u l=1u
M12785 net3805 n4772 net3806 VSS nmos w=1u l=1u
M12786 net3805 n4773 VDD VDD pmos w=2u l=1u
M12787 net3805 n4772 VDD VDD pmos w=2u l=1u
M12788 n4760 net3805 VDD VDD pmos w=2u l=1u
M12789 n4753 net3807 VSS VSS nmos w=1u l=1u
M12790 net3808 n4750 VSS VSS nmos w=1u l=1u
M12791 net3807 n4751 net3808 VSS nmos w=1u l=1u
M12792 net3807 n4750 VDD VDD pmos w=2u l=1u
M12793 net3807 n4751 VDD VDD pmos w=2u l=1u
M12794 n4753 net3807 VDD VDD pmos w=2u l=1u
M12795 N2223 n4774 net3809 VSS nmos w=1u l=1u
M12796 net3809 n4750 VSS VSS nmos w=1u l=1u
M12797 N2223 n4774 VDD VDD pmos w=2u l=1u
M12798 N2223 n4750 VDD VDD pmos w=2u l=1u
M12799 n4774 N1 net3810 VSS nmos w=1u l=1u
M12800 net3810 n4775 VSS VSS nmos w=1u l=1u
M12801 n4774 N1 VDD VDD pmos w=2u l=1u
M12802 n4774 n4775 VDD VDD pmos w=2u l=1u
M12803 n4775 n3257 VSS VSS nmos w=1u l=1u
M12804 n4775 n4776 VSS VSS nmos w=1u l=1u
M12805 n4775 n3257 net3811 VDD pmos w=2u l=1u
M12806 net3811 n4776 VDD VDD pmos w=2u l=1u
M12807 n3257 N324 VDD VDD pmos w=2u l=1u
M12808 n3257 N324 VSS VSS nmos w=1u l=1u
M12809 n4750 n4777 net3812 VSS nmos w=1u l=1u
M12810 net3812 n4776 VSS VSS nmos w=1u l=1u
M12811 n4750 n4777 VDD VDD pmos w=2u l=1u
M12812 n4750 n4776 VDD VDD pmos w=2u l=1u
M12813 n4777 N324 net3813 VSS nmos w=1u l=1u
M12814 net3813 N1 VSS VSS nmos w=1u l=1u
M12815 n4777 N324 VDD VDD pmos w=2u l=1u
M12816 n4777 N1 VDD VDD pmos w=2u l=1u
M12817 n4776 net3814 VSS VSS nmos w=1u l=1u
M12818 net3815 n4778 VSS VSS nmos w=1u l=1u
M12819 net3814 n4751 net3815 VSS nmos w=1u l=1u
M12820 net3814 n4778 VDD VDD pmos w=2u l=1u
M12821 net3814 n4751 VDD VDD pmos w=2u l=1u
M12822 n4776 net3814 VDD VDD pmos w=2u l=1u
M12823 n4778 n4780 net3816 VSS nmos w=1u l=1u
M12824 net3816 n4779 VSS VSS nmos w=1u l=1u
M12825 n4778 n4780 VDD VDD pmos w=2u l=1u
M12826 n4778 n4779 VDD VDD pmos w=2u l=1u
M12827 n4751 net3817 VSS VSS nmos w=1u l=1u
M12828 net3817 n4780 VSS VSS nmos w=1u l=1u
M12829 net3817 n4779 VSS VSS nmos w=1u l=1u
M12830 net3817 n4779 net3818 VDD pmos w=2u l=1u
M12831 n4751 net3817 VDD VDD pmos w=2u l=1u
M12832 net3818 n4780 VDD VDD pmos w=2u l=1u
M12833 n4779 net3819 VSS VSS nmos w=1u l=1u
M12834 net3820 n4782 VSS VSS nmos w=1u l=1u
M12835 net3819 n4781 net3820 VSS nmos w=1u l=1u
M12836 net3819 n4782 VDD VDD pmos w=2u l=1u
M12837 net3819 n4781 VDD VDD pmos w=2u l=1u
M12838 n4779 net3819 VDD VDD pmos w=2u l=1u
M12839 n4780 n4783 net3821 VSS nmos w=1u l=1u
M12840 net3821 n4772 VSS VSS nmos w=1u l=1u
M12841 n4780 n4783 VDD VDD pmos w=2u l=1u
M12842 n4780 n4772 VDD VDD pmos w=2u l=1u
M12843 n4783 N18 net3822 VSS nmos w=1u l=1u
M12844 net3822 n4784 VSS VSS nmos w=1u l=1u
M12845 n4783 N18 VDD VDD pmos w=2u l=1u
M12846 n4783 n4784 VDD VDD pmos w=2u l=1u
M12847 n4784 n3411 VSS VSS nmos w=1u l=1u
M12848 n4784 n4785 VSS VSS nmos w=1u l=1u
M12849 n4784 n3411 net3823 VDD pmos w=2u l=1u
M12850 net3823 n4785 VDD VDD pmos w=2u l=1u
M12851 n4772 n4786 net3824 VSS nmos w=1u l=1u
M12852 net3824 n4785 VSS VSS nmos w=1u l=1u
M12853 n4772 n4786 VDD VDD pmos w=2u l=1u
M12854 n4772 n4785 VDD VDD pmos w=2u l=1u
M12855 n4786 N307 net3825 VSS nmos w=1u l=1u
M12856 net3825 N18 VSS VSS nmos w=1u l=1u
M12857 n4786 N307 VDD VDD pmos w=2u l=1u
M12858 n4786 N18 VDD VDD pmos w=2u l=1u
M12859 n4785 net3826 VSS VSS nmos w=1u l=1u
M12860 net3827 n4787 VSS VSS nmos w=1u l=1u
M12861 net3826 n4773 net3827 VSS nmos w=1u l=1u
M12862 net3826 n4787 VDD VDD pmos w=2u l=1u
M12863 net3826 n4773 VDD VDD pmos w=2u l=1u
M12864 n4785 net3826 VDD VDD pmos w=2u l=1u
M12865 n4787 n4766 net3828 VSS nmos w=1u l=1u
M12866 net3828 n4788 VSS VSS nmos w=1u l=1u
M12867 n4787 n4766 VDD VDD pmos w=2u l=1u
M12868 n4787 n4788 VDD VDD pmos w=2u l=1u
M12869 n4788 n4789 VDD VDD pmos w=2u l=1u
M12870 n4788 n4789 VSS VSS nmos w=1u l=1u
M12871 n4773 n4790 net3829 VSS nmos w=1u l=1u
M12872 net3829 n4789 VSS VSS nmos w=1u l=1u
M12873 n4773 n4790 VDD VDD pmos w=2u l=1u
M12874 n4773 n4789 VDD VDD pmos w=2u l=1u
M12875 n4790 n4766 net3830 VSS nmos w=1u l=1u
M12876 net3830 n4791 VSS VSS nmos w=1u l=1u
M12877 n4790 n4766 VDD VDD pmos w=2u l=1u
M12878 n4790 n4791 VDD VDD pmos w=2u l=1u
M12879 n4766 N52 net3831 VSS nmos w=1u l=1u
M12880 net3831 n4792 VSS VSS nmos w=1u l=1u
M12881 n4766 N52 VDD VDD pmos w=2u l=1u
M12882 n4766 n4792 VDD VDD pmos w=2u l=1u
M12883 n4791 n4794 net3832 VSS nmos w=1u l=1u
M12884 net3832 n4793 VSS VSS nmos w=1u l=1u
M12885 n4791 n4794 VDD VDD pmos w=2u l=1u
M12886 n4791 n4793 VDD VDD pmos w=2u l=1u
M12887 n4794 N273 net3833 VSS nmos w=1u l=1u
M12888 net3833 N52 VSS VSS nmos w=1u l=1u
M12889 n4794 N273 VDD VDD pmos w=2u l=1u
M12890 n4794 N52 VDD VDD pmos w=2u l=1u
M12891 n4793 N290 net3834 VSS nmos w=1u l=1u
M12892 net3834 N35 VSS VSS nmos w=1u l=1u
M12893 n4793 N290 VDD VDD pmos w=2u l=1u
M12894 n4793 N35 VDD VDD pmos w=2u l=1u
M12895 N1901 n4795 net3835 VSS nmos w=1u l=1u
M12896 net3835 n4782 VSS VSS nmos w=1u l=1u
M12897 N1901 n4795 VDD VDD pmos w=2u l=1u
M12898 N1901 n4782 VDD VDD pmos w=2u l=1u
M12899 n4795 N1 net3836 VSS nmos w=1u l=1u
M12900 net3836 n4796 VSS VSS nmos w=1u l=1u
M12901 n4795 N1 VDD VDD pmos w=2u l=1u
M12902 n4795 n4796 VDD VDD pmos w=2u l=1u
M12903 n4796 n3411 VSS VSS nmos w=1u l=1u
M12904 n4796 n4797 VSS VSS nmos w=1u l=1u
M12905 n4796 n3411 net3837 VDD pmos w=2u l=1u
M12906 net3837 n4797 VDD VDD pmos w=2u l=1u
M12907 n3411 N307 VDD VDD pmos w=2u l=1u
M12908 n3411 N307 VSS VSS nmos w=1u l=1u
M12909 n4782 n4798 net3838 VSS nmos w=1u l=1u
M12910 net3838 n4797 VSS VSS nmos w=1u l=1u
M12911 n4782 n4798 VDD VDD pmos w=2u l=1u
M12912 n4782 n4797 VDD VDD pmos w=2u l=1u
M12913 n4798 N307 net3839 VSS nmos w=1u l=1u
M12914 net3839 N1 VSS VSS nmos w=1u l=1u
M12915 n4798 N307 VDD VDD pmos w=2u l=1u
M12916 n4798 N1 VDD VDD pmos w=2u l=1u
M12917 n4797 net3840 VSS VSS nmos w=1u l=1u
M12918 net3841 n4799 VSS VSS nmos w=1u l=1u
M12919 net3840 n4781 net3841 VSS nmos w=1u l=1u
M12920 net3840 n4799 VDD VDD pmos w=2u l=1u
M12921 net3840 n4781 VDD VDD pmos w=2u l=1u
M12922 n4797 net3840 VDD VDD pmos w=2u l=1u
M12923 n4799 n4789 net3842 VSS nmos w=1u l=1u
M12924 net3842 n4800 VSS VSS nmos w=1u l=1u
M12925 n4799 n4789 VDD VDD pmos w=2u l=1u
M12926 n4799 n4800 VDD VDD pmos w=2u l=1u
M12927 n4781 n4802 net3843 VSS nmos w=1u l=1u
M12928 net3843 n4801 VSS VSS nmos w=1u l=1u
M12929 n4781 n4802 VDD VDD pmos w=2u l=1u
M12930 n4781 n4801 VDD VDD pmos w=2u l=1u
M12931 n4802 n4789 net3844 VSS nmos w=1u l=1u
M12932 net3844 n4803 VSS VSS nmos w=1u l=1u
M12933 n4802 n4789 VDD VDD pmos w=2u l=1u
M12934 n4802 n4803 VDD VDD pmos w=2u l=1u
M12935 n4789 N18 net3845 VSS nmos w=1u l=1u
M12936 net3845 n4792 VSS VSS nmos w=1u l=1u
M12937 n4789 N18 VDD VDD pmos w=2u l=1u
M12938 n4789 n4792 VDD VDD pmos w=2u l=1u
M12939 n4792 n3456 VSS VSS nmos w=1u l=1u
M12940 n4792 n3898 VSS VSS nmos w=1u l=1u
M12941 n4792 n3456 net3846 VDD pmos w=2u l=1u
M12942 net3846 n3898 VDD VDD pmos w=2u l=1u
M12943 n3456 N35 VDD VDD pmos w=2u l=1u
M12944 n3456 N35 VSS VSS nmos w=1u l=1u
M12945 n3898 n3741 VDD VDD pmos w=2u l=1u
M12946 n3898 n3741 VSS VSS nmos w=1u l=1u
M12947 n3741 n3745 VSS VSS nmos w=1u l=1u
M12948 n3741 n3746 VSS VSS nmos w=1u l=1u
M12949 n3741 n3745 net3847 VDD pmos w=2u l=1u
M12950 net3847 n3746 VDD VDD pmos w=2u l=1u
M12951 n4803 n4805 net3848 VSS nmos w=1u l=1u
M12952 net3848 n4804 VSS VSS nmos w=1u l=1u
M12953 n4803 n4805 VDD VDD pmos w=2u l=1u
M12954 n4803 n4804 VDD VDD pmos w=2u l=1u
M12955 n4805 N273 net3849 VSS nmos w=1u l=1u
M12956 net3849 N35 VSS VSS nmos w=1u l=1u
M12957 n4805 N273 VDD VDD pmos w=2u l=1u
M12958 n4805 N35 VDD VDD pmos w=2u l=1u
M12959 n4804 N290 net3850 VSS nmos w=1u l=1u
M12960 net3850 N18 VSS VSS nmos w=1u l=1u
M12961 n4804 N290 VDD VDD pmos w=2u l=1u
M12962 n4804 N18 VDD VDD pmos w=2u l=1u
M12963 N1581 n4806 VSS VSS nmos w=1u l=1u
M12964 N1581 n4800 VSS VSS nmos w=1u l=1u
M12965 N1581 n4806 net3851 VDD pmos w=2u l=1u
M12966 net3851 n4800 VDD VDD pmos w=2u l=1u
M12967 n4806 n4808 VSS VSS nmos w=1u l=1u
M12968 n4806 n4807 VSS VSS nmos w=1u l=1u
M12969 n4806 n4808 net3852 VDD pmos w=2u l=1u
M12970 net3852 n4807 VDD VDD pmos w=2u l=1u
M12971 n4808 net3853 VSS VSS nmos w=1u l=1u
M12972 net3854 N1 VSS VSS nmos w=1u l=1u
M12973 net3853 N290 net3854 VSS nmos w=1u l=1u
M12974 net3853 N1 VDD VDD pmos w=2u l=1u
M12975 net3853 N290 VDD VDD pmos w=2u l=1u
M12976 n4808 net3853 VDD VDD pmos w=2u l=1u
M12977 n4807 n3603 VSS VSS nmos w=1u l=1u
M12978 n4807 n3746 VSS VSS nmos w=1u l=1u
M12979 n4807 n3603 net3855 VDD pmos w=2u l=1u
M12980 net3855 n3746 VDD VDD pmos w=2u l=1u
M12981 n4800 n4801 VDD VDD pmos w=2u l=1u
M12982 n4800 n4801 VSS VSS nmos w=1u l=1u
M12983 n4801 N545 net3856 VSS nmos w=1u l=1u
M12984 net3856 n4809 VSS VSS nmos w=1u l=1u
M12985 n4801 N545 VDD VDD pmos w=2u l=1u
M12986 n4801 n4809 VDD VDD pmos w=2u l=1u
M12987 N545 n3746 VSS VSS nmos w=1u l=1u
M12988 N545 n3929 VSS VSS nmos w=1u l=1u
M12989 N545 n3746 net3857 VDD pmos w=2u l=1u
M12990 net3857 n3929 VDD VDD pmos w=2u l=1u
M12991 n3929 N1 VDD VDD pmos w=2u l=1u
M12992 n3929 N1 VSS VSS nmos w=1u l=1u
M12993 n4809 n3603 VSS VSS nmos w=1u l=1u
M12994 n4809 n3745 VSS VSS nmos w=1u l=1u
M12995 n4809 n3603 net3858 VDD pmos w=2u l=1u
M12996 net3858 n3745 VDD VDD pmos w=2u l=1u
M12997 n3603 N18 VDD VDD pmos w=2u l=1u
M12998 n3603 N18 VSS VSS nmos w=1u l=1u
M12999 n3745 N290 VSS VSS nmos w=1u l=1u
M13000 n3745 n3746 VSS VSS nmos w=1u l=1u
M13001 n3745 N290 net3859 VDD pmos w=2u l=1u
M13002 net3859 n3746 VDD VDD pmos w=2u l=1u
M13003 n3746 N273 VDD VDD pmos w=2u l=1u
M13004 n3746 N273 VSS VSS nmos w=1u l=1u
.ENDS

